--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/

-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC
-- Version: 2013.4
-- Copyright (C) 2013 Xilinx Inc. All rights reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity huffman_decoder is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    code_V_V_dout : IN STD_LOGIC_VECTOR (31 downto 0);
    code_V_V_empty_n : IN STD_LOGIC;
    code_V_V_read : OUT STD_LOGIC;
    z1_V_V_din : OUT STD_LOGIC_VECTOR (13 downto 0);
    z1_V_V_full_n : IN STD_LOGIC;
    z1_V_V_write : OUT STD_LOGIC;
    z2_V_V_din : OUT STD_LOGIC_VECTOR (2 downto 0);
    z2_V_V_full_n : IN STD_LOGIC;
    z2_V_V_write : OUT STD_LOGIC;
    ap_return : OUT STD_LOGIC_VECTOR (0 downto 0) );
end;


architecture behav of huffman_decoder is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "huffman_decoder,hls_ip_2013_4,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020clg484-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.664000,HLS_SYN_LAT=67841,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=0,HLS_SYN_LUT=0}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_st1_fsm_0 : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    constant ap_ST_st2_fsm_1 : STD_LOGIC_VECTOR (3 downto 0) := "0001";
    constant ap_ST_st3_fsm_2 : STD_LOGIC_VECTOR (3 downto 0) := "0010";
    constant ap_ST_st4_fsm_3 : STD_LOGIC_VECTOR (3 downto 0) := "0011";
    constant ap_ST_st5_fsm_4 : STD_LOGIC_VECTOR (3 downto 0) := "0100";
    constant ap_ST_st6_fsm_5 : STD_LOGIC_VECTOR (3 downto 0) := "0101";
    constant ap_ST_st7_fsm_6 : STD_LOGIC_VECTOR (3 downto 0) := "0110";
    constant ap_ST_st8_fsm_7 : STD_LOGIC_VECTOR (3 downto 0) := "0111";
    constant ap_ST_st9_fsm_8 : STD_LOGIC_VECTOR (3 downto 0) := "1000";
    constant ap_ST_st10_fsm_9 : STD_LOGIC_VECTOR (3 downto 0) := "1001";
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv96_0 : STD_LOGIC_VECTOR (95 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv7_0 : STD_LOGIC_VECTOR (6 downto 0) := "0000000";
    constant ap_const_lv9_0 : STD_LOGIC_VECTOR (8 downto 0) := "000000000";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_lv9_100 : STD_LOGIC_VECTOR (8 downto 0) := "100000000";
    constant ap_const_lv9_1 : STD_LOGIC_VECTOR (8 downto 0) := "000000001";
    constant ap_const_lv7_41 : STD_LOGIC_VECTOR (6 downto 0) := "1000001";
    constant ap_const_lv7_20 : STD_LOGIC_VECTOR (6 downto 0) := "0100000";
    constant ap_const_lv32_10 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010000";
    constant ap_const_lv32_22 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000100010";
    constant ap_const_lv32_6 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000110";
    constant ap_const_lv7_1 : STD_LOGIC_VECTOR (6 downto 0) := "0000001";
    constant ap_const_lv32_1 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000001";
    constant ap_const_lv19_7FFFF : STD_LOGIC_VECTOR (18 downto 0) := "1111111111111111111";
    constant ap_const_lv32_4 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000100";
    constant ap_const_lv32_5 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000101";
    constant ap_const_lv32_2 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000010";
    constant ap_const_lv32_3 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000011";
    constant ap_const_lv10_10 : STD_LOGIC_VECTOR (9 downto 0) := "0000010000";
    constant ap_const_lv32_9 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001001";
    constant ap_const_lv10_3F0 : STD_LOGIC_VECTOR (9 downto 0) := "1111110000";
    constant ap_const_lv10_0 : STD_LOGIC_VECTOR (9 downto 0) := "0000000000";
    constant ap_const_lv32_1F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011111";
    constant ap_const_lv7_70 : STD_LOGIC_VECTOR (6 downto 0) := "1110000";
    constant ap_const_lv32_8 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001000";
    constant ap_const_lv32_F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001111";
    constant ap_const_lv11_0 : STD_LOGIC_VECTOR (10 downto 0) := "00000000000";
    constant ap_const_lv1_1 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv2_1 : STD_LOGIC_VECTOR (1 downto 0) := "01";
    constant ap_const_lv2_2 : STD_LOGIC_VECTOR (1 downto 0) := "10";
    constant ap_const_lv2_0 : STD_LOGIC_VECTOR (1 downto 0) := "00";
    constant ap_const_lv3_1 : STD_LOGIC_VECTOR (2 downto 0) := "001";

    signal ap_CS_fsm : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal val_table_address0 : STD_LOGIC_VECTOR (5 downto 0);
    signal val_table_ce0 : STD_LOGIC;
    signal val_table_q0 : STD_LOGIC_VECTOR (5 downto 0);
    signal bit_cnt_table_address0 : STD_LOGIC_VECTOR (5 downto 0);
    signal bit_cnt_table_ce0 : STD_LOGIC;
    signal bit_cnt_table_q0 : STD_LOGIC_VECTOR (4 downto 0);
    signal dec_e_table_address0 : STD_LOGIC_VECTOR (5 downto 0);
    signal dec_e_table_ce0 : STD_LOGIC;
    signal dec_e_table_q0 : STD_LOGIC_VECTOR (18 downto 0);
    signal tmp_fu_321_p2 : STD_LOGIC_VECTOR (8 downto 0);
    signal tmp_reg_913 : STD_LOGIC_VECTOR (8 downto 0);
    signal r_V_10_fu_347_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_1_fu_327_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_2_nbreadreq_fu_134_p3 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_sig_bdd_76 : BOOLEAN;
    signal data_reg_count_V_fu_353_p2 : STD_LOGIC_VECTOR (6 downto 0);
    signal full_e_V_reg_934 : STD_LOGIC_VECTOR (18 downto 0);
    signal inner_cnt_4_cast_fu_369_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal inner_cnt_4_cast_reg_939 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_4_fu_373_p3 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_4_reg_945 : STD_LOGIC_VECTOR (0 downto 0);
    signal j_fu_381_p2 : STD_LOGIC_VECTOR (6 downto 0);
    signal j_reg_949 : STD_LOGIC_VECTOR (6 downto 0);
    signal dec_e_table_load_reg_969 : STD_LOGIC_VECTOR (18 downto 0);
    signal bt_cnt_V_reg_974 : STD_LOGIC_VECTOR (4 downto 0);
    signal tmp_s_fu_422_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_12_reg_988 : STD_LOGIC_VECTOR (1 downto 0);
    signal zh_2_1_V_reg_993 : STD_LOGIC_VECTOR (0 downto 0);
    signal zh_2_2_V_fu_471_p1 : STD_LOGIC_VECTOR (0 downto 0);
    signal zh_2_2_V_reg_1002 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_13_fu_479_p3 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_13_reg_1010 : STD_LOGIC_VECTOR (9 downto 0);
    signal op2_assign_fu_491_p2 : STD_LOGIC_VECTOR (9 downto 0);
    signal op2_assign_reg_1015 : STD_LOGIC_VECTOR (9 downto 0);
    signal signs_V_fu_547_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal signs_V_reg_1020 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_35_fu_551_p1 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_35_reg_1025 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_21_fu_555_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_21_reg_1030 : STD_LOGIC_VECTOR (0 downto 0);
    signal r_V_s_reg_1038 : STD_LOGIC_VECTOR (30 downto 0);
    signal p_neg1_fu_581_p2 : STD_LOGIC_VECTOR (6 downto 0);
    signal p_neg1_reg_1043 : STD_LOGIC_VECTOR (6 downto 0);
    signal tmp_V_2_fu_702_p3 : STD_LOGIC_VECTOR (10 downto 0);
    signal tmp_V_2_reg_1048 : STD_LOGIC_VECTOR (10 downto 0);
    signal ap_sig_bdd_142 : BOOLEAN;
    signal tmp_38_fu_780_p1 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_38_reg_1053 : STD_LOGIC_VECTOR (0 downto 0);
    signal p_0554_3_fu_801_p3 : STD_LOGIC_VECTOR (2 downto 0);
    signal p_0554_3_reg_1058 : STD_LOGIC_VECTOR (2 downto 0);
    signal data_reg_count_V_1_fu_840_p2 : STD_LOGIC_VECTOR (6 downto 0);
    signal r_V_14_fu_895_p3 : STD_LOGIC_VECTOR (95 downto 0);
    signal p_s_reg_206 : STD_LOGIC_VECTOR (95 downto 0);
    signal p_1_reg_218 : STD_LOGIC_VECTOR (6 downto 0);
    signal cnt_reg_230 : STD_LOGIC_VECTOR (8 downto 0);
    signal inner_cnt_reg_241 : STD_LOGIC_VECTOR (31 downto 0);
    signal inner_cnt_3_reg_297 : STD_LOGIC_VECTOR (31 downto 0);
    signal lhs_V_reg_253 : STD_LOGIC_VECTOR (95 downto 0);
    signal exitcond_fu_315_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal p_0622_1_reg_264 : STD_LOGIC_VECTOR (6 downto 0);
    signal inner_cnt_2_reg_275 : STD_LOGIC_VECTOR (6 downto 0);
    signal inner_cnt_1_reg_286 : STD_LOGIC_VECTOR (31 downto 0);
    signal inner_cnt_3_phi_fu_301_p4 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_5_fu_387_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal tmp_6_fu_393_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal tmp_10_fu_435_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal inner_cnt_3_phi_fu_301_p4_temp: signed (32-1 downto 0);
    signal tmp_V_6_cast_fu_637_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal tmp_V_1_fu_630_p3_temp: signed (11-1 downto 0);
    signal tmp_V_7_cast_fu_811_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal tmp_V_2_reg_1048_temp: signed (11-1 downto 0);
    signal tmp_V_4_fu_768_p1 : STD_LOGIC_VECTOR (2 downto 0);
    signal tmp_V_3_fu_761_p3_temp: signed (2-1 downto 0);
    signal tmp_V_5_fu_832_p1 : STD_LOGIC_VECTOR (2 downto 0);
    signal tmp_V_6_fu_825_p3_temp: signed (2-1 downto 0);
    signal e_length_V_1_fu_130 : STD_LOGIC_VECTOR (8 downto 0);
    signal e_length_V_fu_427_p1 : STD_LOGIC_VECTOR (8 downto 0);
    signal temp_V_fu_333_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_7_fu_337_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal r_V_9_fu_341_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_8_fu_398_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_9_fu_401_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal tmp_16_fu_407_p1 : STD_LOGIC_VECTOR (18 downto 0);
    signal tmp_11_cast_fu_411_p2 : STD_LOGIC_VECTOR (18 downto 0);
    signal tmp_3_fu_417_p2 : STD_LOGIC_VECTOR (18 downto 0);
    signal tmp_11_fu_443_p4 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_32_fu_475_p1 : STD_LOGIC_VECTOR (7 downto 0);
    signal op2_assign_fu_491_p0 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_23_cast_fu_487_p1 : STD_LOGIC_VECTOR (9 downto 0);
    signal e_length_V_1_fu_130_temp: signed (9-1 downto 0);
    signal tmp_15_fu_509_p0 : STD_LOGIC_VECTOR (63 downto 0);
    signal op2_assign_fu_491_p2_temp: signed (10-1 downto 0);
    signal tmp_15_fu_509_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_18_fu_519_p1 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_18_fu_519_p2 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_19_fu_529_p0 : STD_LOGIC_VECTOR (63 downto 0);
    signal tmp_18_fu_519_p2_temp: signed (10-1 downto 0);
    signal tmp_19_fu_529_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_33_fu_501_p3 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_20_fu_533_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_17_fu_513_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal r_V_fu_539_p3 : STD_LOGIC_VECTOR (95 downto 0);
    signal p_neg_fu_575_p2 : STD_LOGIC_VECTOR (6 downto 0);
    signal tmp_39_fu_571_p1 : STD_LOGIC_VECTOR (6 downto 0);
    signal phitmp_fu_590_p4 : STD_LOGIC_VECTOR (7 downto 0);
    signal tmp_14_fu_603_p3 : STD_LOGIC_VECTOR (9 downto 0);
    signal z1_1_V_cast_fu_600_p1 : STD_LOGIC_VECTOR (10 downto 0);
    signal z1_1_V_fu_614_p2 : STD_LOGIC_VECTOR (10 downto 0);
    signal p_s_16_fu_620_p3 : STD_LOGIC_VECTOR (10 downto 0);
    signal tmp_V_1_fu_630_p3 : STD_LOGIC_VECTOR (10 downto 0);
    signal r_V_11_fu_627_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal signs_V_2_fu_642_p3 : STD_LOGIC_VECTOR (31 downto 0);
    signal not_tmp_s_fu_652_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal z1_2_V_cast_fu_610_p1 : STD_LOGIC_VECTOR (10 downto 0);
    signal tmp_36_fu_648_p1 : STD_LOGIC_VECTOR (0 downto 0);
    signal z1_2_V_fu_667_p2 : STD_LOGIC_VECTOR (10 downto 0);
    signal r_V_1_fu_681_p4 : STD_LOGIC_VECTOR (30 downto 0);
    signal tmp_22_fu_661_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal p_1_17_fu_673_p3 : STD_LOGIC_VECTOR (10 downto 0);
    signal r_V_12_fu_691_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal signs_V_4_fu_710_p3 : STD_LOGIC_VECTOR (31 downto 0);
    signal p_5_cast_fu_657_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal sign_cnt_V_fu_695_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_37_fu_718_p1 : STD_LOGIC_VECTOR (0 downto 0);
    signal phitmp1761_s_fu_733_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal zh_2_1_V_reg_993_temp: signed (1-1 downto 0);
    signal zh_2_1_V_cast_fu_587_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal r_V_2_fu_741_p4 : STD_LOGIC_VECTOR (30 downto 0);
    signal p_0554_1_fu_722_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal phitmp1761_s_fu_733_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_V_3_fu_761_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal r_V_13_fu_751_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal signs_V_6_fu_773_p3 : STD_LOGIC_VECTOR (31 downto 0);
    signal sign_cnt_V_1_fu_755_p2 : STD_LOGIC_VECTOR (1 downto 0);
    signal p_0554_2_fu_784_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal p_0554_2_cast_fu_791_p1 : STD_LOGIC_VECTOR (2 downto 0);
    signal sign_cnt_V_2_fu_795_p2 : STD_LOGIC_VECTOR (2 downto 0);
    signal phitmp1763_s_fu_818_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal zh_2_2_V_reg_1002_temp: signed (1-1 downto 0);
    signal zh_2_2_V_cast_fu_808_p1 : STD_LOGIC_VECTOR (1 downto 0);
    signal phitmp1763_s_fu_818_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_V_6_fu_825_p3 : STD_LOGIC_VECTOR (1 downto 0);
    signal tmp_23_fu_837_p1 : STD_LOGIC_VECTOR (6 downto 0);
    signal tmp_44_cast_fu_845_p1 : STD_LOGIC_VECTOR (9 downto 0);
    signal op2_assign_1_fu_848_p2 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_24_fu_865_p0 : STD_LOGIC_VECTOR (63 downto 0);
    signal op2_assign_1_fu_848_p2_temp: signed (10-1 downto 0);
    signal tmp_24_fu_865_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_26_fu_875_p2 : STD_LOGIC_VECTOR (9 downto 0);
    signal tmp_27_fu_885_p0 : STD_LOGIC_VECTOR (63 downto 0);
    signal tmp_26_fu_875_p2_temp: signed (10-1 downto 0);
    signal tmp_27_fu_885_p1 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_40_fu_857_p3 : STD_LOGIC_VECTOR (0 downto 0);
    signal tmp_28_fu_889_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal tmp_25_fu_869_p2 : STD_LOGIC_VECTOR (95 downto 0);
    signal ap_NS_fsm : STD_LOGIC_VECTOR (3 downto 0);

    component huffman_decoder_val_table IS
    generic (
        DataWidth : INTEGER;
        AddressRange : INTEGER;
        AddressWidth : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        address0 : IN STD_LOGIC_VECTOR (5 downto 0);
        ce0 : IN STD_LOGIC;
        q0 : OUT STD_LOGIC_VECTOR (5 downto 0) );
    end component;


    component huffman_decoder_bit_cnt_table IS
    generic (
        DataWidth : INTEGER;
        AddressRange : INTEGER;
        AddressWidth : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        address0 : IN STD_LOGIC_VECTOR (5 downto 0);
        ce0 : IN STD_LOGIC;
        q0 : OUT STD_LOGIC_VECTOR (4 downto 0) );
    end component;


    component huffman_decoder_dec_e_table IS
    generic (
        DataWidth : INTEGER;
        AddressRange : INTEGER;
        AddressWidth : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        address0 : IN STD_LOGIC_VECTOR (5 downto 0);
        ce0 : IN STD_LOGIC;
        q0 : OUT STD_LOGIC_VECTOR (18 downto 0) );
    end component;



begin
    val_table_U : component huffman_decoder_val_table
    generic map (
        DataWidth => 6,
        AddressRange => 64,
        AddressWidth => 6)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        address0 => val_table_address0,
        ce0 => val_table_ce0,
        q0 => val_table_q0);

    bit_cnt_table_U : component huffman_decoder_bit_cnt_table
    generic map (
        DataWidth => 5,
        AddressRange => 64,
        AddressWidth => 6)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        address0 => bit_cnt_table_address0,
        ce0 => bit_cnt_table_ce0,
        q0 => bit_cnt_table_q0);

    dec_e_table_U : component huffman_decoder_dec_e_table
    generic map (
        DataWidth => 19,
        AddressRange => 64,
        AddressWidth => 6)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        address0 => dec_e_table_address0,
        ce0 => dec_e_table_ce0,
        q0 => dec_e_table_q0);





    -- the current state (ap_CS_fsm) of the state machine. --
    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_CS_fsm <= ap_ST_st1_fsm_0;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    -- cnt_reg_230 assign process. --
    cnt_reg_230_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm))) then 
                cnt_reg_230 <= tmp_reg_913;
            elsif (((ap_ST_st1_fsm_0 = ap_CS_fsm) and not((ap_start = ap_const_logic_0)))) then 
                cnt_reg_230 <= ap_const_lv9_0;
            end if; 
        end if;
    end process;

    -- e_length_V_1_fu_130 assign process. --
    e_length_V_1_fu_130_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st7_fsm_6 = ap_CS_fsm) and (ap_const_lv1_0 = tmp_4_reg_945) and not((ap_const_lv1_0 = tmp_s_fu_422_p2)))) then 
                e_length_V_1_fu_130(0) <= e_length_V_fu_427_p1(0);
                e_length_V_1_fu_130(1) <= e_length_V_fu_427_p1(1);
                e_length_V_1_fu_130(2) <= e_length_V_fu_427_p1(2);
                e_length_V_1_fu_130(3) <= e_length_V_fu_427_p1(3);
                e_length_V_1_fu_130(4) <= e_length_V_fu_427_p1(4);
            elsif (((ap_ST_st1_fsm_0 = ap_CS_fsm) and not((ap_start = ap_const_logic_0)))) then 
                e_length_V_1_fu_130(0) <= '0';
                e_length_V_1_fu_130(1) <= '0';
                e_length_V_1_fu_130(2) <= '0';
                e_length_V_1_fu_130(3) <= '0';
                e_length_V_1_fu_130(4) <= '0';
            end if; 
        end if;
    end process;

    -- inner_cnt_1_reg_286 assign process. --
    inner_cnt_1_reg_286_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st7_fsm_6 = ap_CS_fsm) and (ap_const_lv1_0 = tmp_4_reg_945) and (ap_const_lv1_0 = tmp_s_fu_422_p2))) then 
                inner_cnt_1_reg_286 <= inner_cnt_4_cast_reg_939;
            elsif (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not(ap_sig_bdd_76) and ((tmp_1_fu_327_p2 = ap_const_lv1_0) or (ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)))) then 
                inner_cnt_1_reg_286 <= inner_cnt_reg_241;
            end if; 
        end if;
    end process;

    -- inner_cnt_2_reg_275 assign process. --
    inner_cnt_2_reg_275_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st7_fsm_6 = ap_CS_fsm) and (ap_const_lv1_0 = tmp_4_reg_945) and (ap_const_lv1_0 = tmp_s_fu_422_p2))) then 
                inner_cnt_2_reg_275 <= j_reg_949;
            elsif (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not(ap_sig_bdd_76) and ((tmp_1_fu_327_p2 = ap_const_lv1_0) or (ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)))) then 
                inner_cnt_2_reg_275 <= ap_const_lv7_0;
            end if; 
        end if;
    end process;

    -- inner_cnt_3_reg_297 assign process. --
    inner_cnt_3_reg_297_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st4_fsm_3 = ap_CS_fsm) and not((ap_const_lv1_0 = tmp_4_fu_373_p3)))) then 
                inner_cnt_3_reg_297 <= inner_cnt_1_reg_286;
            elsif (((ap_ST_st7_fsm_6 = ap_CS_fsm) and (ap_const_lv1_0 = tmp_4_reg_945) and not((ap_const_lv1_0 = tmp_s_fu_422_p2)))) then 
                inner_cnt_3_reg_297 <= inner_cnt_4_cast_reg_939;
            end if; 
        end if;
    end process;

    -- inner_cnt_reg_241 assign process. --
    inner_cnt_reg_241_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm))) then 
                inner_cnt_reg_241 <= inner_cnt_3_reg_297;
            elsif (((ap_ST_st1_fsm_0 = ap_CS_fsm) and not((ap_start = ap_const_logic_0)))) then 
                inner_cnt_reg_241 <= ap_const_lv32_0;
            end if; 
        end if;
    end process;

    -- lhs_V_reg_253 assign process. --
    lhs_V_reg_253_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st2_fsm_1 = ap_CS_fsm) and (ap_const_lv1_0 = exitcond_fu_315_p2))) then 
                lhs_V_reg_253 <= p_s_reg_206;
            elsif (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not((tmp_1_fu_327_p2 = ap_const_lv1_0)) and not((ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)) and not(ap_sig_bdd_76))) then 
                lhs_V_reg_253 <= r_V_10_fu_347_p2;
            end if; 
        end if;
    end process;

    -- p_0622_1_reg_264 assign process. --
    p_0622_1_reg_264_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st2_fsm_1 = ap_CS_fsm) and (ap_const_lv1_0 = exitcond_fu_315_p2))) then 
                p_0622_1_reg_264 <= p_1_reg_218;
            elsif (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not((tmp_1_fu_327_p2 = ap_const_lv1_0)) and not((ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)) and not(ap_sig_bdd_76))) then 
                p_0622_1_reg_264 <= data_reg_count_V_fu_353_p2;
            end if; 
        end if;
    end process;

    -- p_1_reg_218 assign process. --
    p_1_reg_218_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm))) then 
                p_1_reg_218 <= data_reg_count_V_1_fu_840_p2;
            elsif (((ap_ST_st1_fsm_0 = ap_CS_fsm) and not((ap_start = ap_const_logic_0)))) then 
                p_1_reg_218 <= ap_const_lv7_0;
            end if; 
        end if;
    end process;

    -- p_s_reg_206 assign process. --
    p_s_reg_206_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm))) then 
                p_s_reg_206 <= r_V_14_fu_895_p3;
            elsif (((ap_ST_st1_fsm_0 = ap_CS_fsm) and not((ap_start = ap_const_logic_0)))) then 
                p_s_reg_206 <= ap_const_lv96_0;
            end if; 
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_ST_st6_fsm_5 = ap_CS_fsm)) then
                bt_cnt_V_reg_974 <= bit_cnt_table_q0;
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_ST_st5_fsm_4 = ap_CS_fsm)) then
                dec_e_table_load_reg_969 <= dec_e_table_q0;
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not(ap_sig_bdd_76) and ((tmp_1_fu_327_p2 = ap_const_lv1_0) or (ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)))) then
                full_e_V_reg_934 <= lhs_V_reg_253(34 downto 16);
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_ST_st4_fsm_3 = ap_CS_fsm)) then
                inner_cnt_4_cast_reg_939(0) <= inner_cnt_4_cast_fu_369_p1(0);
    inner_cnt_4_cast_reg_939(1) <= inner_cnt_4_cast_fu_369_p1(1);
    inner_cnt_4_cast_reg_939(2) <= inner_cnt_4_cast_fu_369_p1(2);
    inner_cnt_4_cast_reg_939(3) <= inner_cnt_4_cast_fu_369_p1(3);
    inner_cnt_4_cast_reg_939(4) <= inner_cnt_4_cast_fu_369_p1(4);
    inner_cnt_4_cast_reg_939(5) <= inner_cnt_4_cast_fu_369_p1(5);
    inner_cnt_4_cast_reg_939(6) <= inner_cnt_4_cast_fu_369_p1(6);
                j_reg_949 <= j_fu_381_p2;
                tmp_4_reg_945 <= inner_cnt_2_reg_275(6 downto 6);
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_ST_st8_fsm_7 = ap_CS_fsm)) then
                op2_assign_reg_1015 <= op2_assign_fu_491_p2;
                p_neg1_reg_1043 <= p_neg1_fu_581_p2;
                r_V_s_reg_1038 <= r_V_fu_539_p3(31 downto 1);
                signs_V_reg_1020 <= signs_V_fu_547_p1;
                tmp_12_reg_988 <= val_table_q0(3 downto 2);
                tmp_13_reg_1010 <= tmp_13_fu_479_p3;
                tmp_21_reg_1030 <= tmp_21_fu_555_p2;
                tmp_35_reg_1025 <= tmp_35_fu_551_p1;
                zh_2_1_V_reg_993 <= val_table_q0(1 downto 1);
                zh_2_2_V_reg_1002 <= zh_2_2_V_fu_471_p1;
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st9_fsm_8 = ap_CS_fsm) and not(ap_sig_bdd_142))) then
                p_0554_3_reg_1058 <= p_0554_3_fu_801_p3;
                tmp_V_2_reg_1048 <= tmp_V_2_fu_702_p3;
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_ST_st9_fsm_8 = ap_CS_fsm) and not(ap_sig_bdd_142) and not((ap_const_lv1_0 = zh_2_2_V_reg_1002)))) then
                tmp_38_reg_1053 <= tmp_38_fu_780_p1;
            end if;
        end if;
    end process;

    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_ST_st2_fsm_1 = ap_CS_fsm)) then
                tmp_reg_913 <= tmp_fu_321_p2;
            end if;
        end if;
    end process;
    inner_cnt_4_cast_reg_939(31 downto 7) <= "0000000000000000000000000";
    e_length_V_1_fu_130(8 downto 5) <= "0000";

    -- the next state (ap_NS_fsm) of the state machine. --
    ap_NS_fsm_assign_proc : process (ap_start , ap_CS_fsm , tmp_1_fu_327_p2 , tmp_2_nbreadreq_fu_134_p3 , ap_sig_bdd_76 , tmp_4_fu_373_p3 , tmp_4_reg_945 , tmp_s_fu_422_p2 , ap_sig_bdd_142 , exitcond_fu_315_p2)
    begin
        case ap_CS_fsm is
            when ap_ST_st1_fsm_0 => 
                if (not((ap_start = ap_const_logic_0))) then
                    ap_NS_fsm <= ap_ST_st2_fsm_1;
                else
                    ap_NS_fsm <= ap_ST_st1_fsm_0;
                end if;
            when ap_ST_st2_fsm_1 => 
                if (not((ap_const_lv1_0 = exitcond_fu_315_p2))) then
                    ap_NS_fsm <= ap_ST_st1_fsm_0;
                else
                    ap_NS_fsm <= ap_ST_st3_fsm_2;
                end if;
            when ap_ST_st3_fsm_2 => 
                if ((not(ap_sig_bdd_76) and ((tmp_1_fu_327_p2 = ap_const_lv1_0) or (ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)))) then
                    ap_NS_fsm <= ap_ST_st4_fsm_3;
                elsif ((not((tmp_1_fu_327_p2 = ap_const_lv1_0)) and not((ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)) and not(ap_sig_bdd_76))) then
                    ap_NS_fsm <= ap_ST_st3_fsm_2;
                else
                    ap_NS_fsm <= ap_ST_st3_fsm_2;
                end if;
            when ap_ST_st4_fsm_3 => 
                if (not((ap_const_lv1_0 = tmp_4_fu_373_p3))) then
                    ap_NS_fsm <= ap_ST_st7_fsm_6;
                else
                    ap_NS_fsm <= ap_ST_st5_fsm_4;
                end if;
            when ap_ST_st5_fsm_4 => 
                ap_NS_fsm <= ap_ST_st6_fsm_5;
            when ap_ST_st6_fsm_5 => 
                ap_NS_fsm <= ap_ST_st7_fsm_6;
            when ap_ST_st7_fsm_6 => 
                if ((not((ap_const_lv1_0 = tmp_4_reg_945)) or not((ap_const_lv1_0 = tmp_s_fu_422_p2)))) then
                    ap_NS_fsm <= ap_ST_st8_fsm_7;
                else
                    ap_NS_fsm <= ap_ST_st4_fsm_3;
                end if;
            when ap_ST_st8_fsm_7 => 
                ap_NS_fsm <= ap_ST_st9_fsm_8;
            when ap_ST_st9_fsm_8 => 
                if (not(ap_sig_bdd_142)) then
                    ap_NS_fsm <= ap_ST_st10_fsm_9;
                else
                    ap_NS_fsm <= ap_ST_st9_fsm_8;
                end if;
            when ap_ST_st10_fsm_9 => 
                if (not(ap_sig_bdd_142)) then
                    ap_NS_fsm <= ap_ST_st2_fsm_1;
                else
                    ap_NS_fsm <= ap_ST_st10_fsm_9;
                end if;
            when others =>  
                ap_NS_fsm <= "XXXX";
        end case;
    end process;

    -- ap_done assign process. --
    ap_done_assign_proc : process(ap_CS_fsm, exitcond_fu_315_p2)
    begin
        if (((ap_ST_st2_fsm_1 = ap_CS_fsm) and not((ap_const_lv1_0 = exitcond_fu_315_p2)))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;


    -- ap_idle assign process. --
    ap_idle_assign_proc : process(ap_start, ap_CS_fsm)
    begin
        if ((not((ap_const_logic_1 = ap_start)) and (ap_ST_st1_fsm_0 = ap_CS_fsm))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    -- ap_ready assign process. --
    ap_ready_assign_proc : process(ap_CS_fsm, exitcond_fu_315_p2)
    begin
        if (((ap_ST_st2_fsm_1 = ap_CS_fsm) and not((ap_const_lv1_0 = exitcond_fu_315_p2)))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;

    ap_return <= ap_const_lv1_1;

    -- ap_sig_bdd_142 assign process. --
    ap_sig_bdd_142_assign_proc : process(z1_V_V_full_n, z2_V_V_full_n)
    begin
                ap_sig_bdd_142 <= ((z1_V_V_full_n = ap_const_logic_0) or (z2_V_V_full_n = ap_const_logic_0));
    end process;


    -- ap_sig_bdd_76 assign process. --
    ap_sig_bdd_76_assign_proc : process(code_V_V_empty_n, tmp_1_fu_327_p2, tmp_2_nbreadreq_fu_134_p3)
    begin
                ap_sig_bdd_76 <= ((code_V_V_empty_n = ap_const_logic_0) and not((tmp_1_fu_327_p2 = ap_const_lv1_0)) and not((ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)));
    end process;

    bit_cnt_table_address0 <= tmp_6_fu_393_p1(6 - 1 downto 0);

    -- bit_cnt_table_ce0 assign process. --
    bit_cnt_table_ce0_assign_proc : process(ap_CS_fsm)
    begin
        if ((ap_ST_st5_fsm_4 = ap_CS_fsm)) then 
            bit_cnt_table_ce0 <= ap_const_logic_1;
        else 
            bit_cnt_table_ce0 <= ap_const_logic_0;
        end if; 
    end process;


    -- code_V_V_read assign process. --
    code_V_V_read_assign_proc : process(ap_CS_fsm, tmp_1_fu_327_p2, tmp_2_nbreadreq_fu_134_p3, ap_sig_bdd_76)
    begin
        if (((ap_ST_st3_fsm_2 = ap_CS_fsm) and not((tmp_1_fu_327_p2 = ap_const_lv1_0)) and not((ap_const_lv1_0 = tmp_2_nbreadreq_fu_134_p3)) and not(ap_sig_bdd_76))) then 
            code_V_V_read <= ap_const_logic_1;
        else 
            code_V_V_read <= ap_const_logic_0;
        end if; 
    end process;

    data_reg_count_V_1_fu_840_p2 <= std_logic_vector(unsigned(p_neg1_reg_1043) - unsigned(tmp_23_fu_837_p1));
    data_reg_count_V_fu_353_p2 <= std_logic_vector(unsigned(p_0622_1_reg_264) + unsigned(ap_const_lv7_20));
    dec_e_table_address0 <= tmp_5_fu_387_p1(6 - 1 downto 0);

    -- dec_e_table_ce0 assign process. --
    dec_e_table_ce0_assign_proc : process(ap_CS_fsm)
    begin
        if ((ap_ST_st4_fsm_3 = ap_CS_fsm)) then 
            dec_e_table_ce0 <= ap_const_logic_1;
        else 
            dec_e_table_ce0 <= ap_const_logic_0;
        end if; 
    end process;

    e_length_V_fu_427_p1 <= std_logic_vector(resize(unsigned(bt_cnt_V_reg_974),9));
    exitcond_fu_315_p2 <= "1" when (cnt_reg_230 = ap_const_lv9_100) else "0";

    -- inner_cnt_3_phi_fu_301_p4 assign process. --
    inner_cnt_3_phi_fu_301_p4_assign_proc : process(ap_CS_fsm, inner_cnt_4_cast_reg_939, tmp_4_reg_945, tmp_s_fu_422_p2, inner_cnt_3_reg_297)
    begin
        if (((ap_ST_st7_fsm_6 = ap_CS_fsm) and (ap_const_lv1_0 = tmp_4_reg_945) and not((ap_const_lv1_0 = tmp_s_fu_422_p2)))) then 
            inner_cnt_3_phi_fu_301_p4 <= inner_cnt_4_cast_reg_939;
        else 
            inner_cnt_3_phi_fu_301_p4 <= inner_cnt_3_reg_297;
        end if; 
    end process;

    inner_cnt_4_cast_fu_369_p1 <= std_logic_vector(resize(unsigned(inner_cnt_2_reg_275),32));
    j_fu_381_p2 <= std_logic_vector(unsigned(inner_cnt_2_reg_275) + unsigned(ap_const_lv7_1));
    not_tmp_s_fu_652_p2 <= (tmp_21_reg_1030 xor ap_const_lv1_1);
    op2_assign_1_fu_848_p2 <= std_logic_vector(unsigned(op2_assign_reg_1015) + unsigned(tmp_44_cast_fu_845_p1));
    op2_assign_fu_491_p0 <= tmp_23_cast_fu_487_p1;
    op2_assign_fu_491_p2 <= std_logic_vector(unsigned(op2_assign_fu_491_p0) + unsigned(ap_const_lv10_10));
    p_0554_1_fu_722_p3 <= 
        p_5_cast_fu_657_p1 when (tmp_22_fu_661_p2(0) = '1') else 
        sign_cnt_V_fu_695_p3;
    p_0554_2_cast_fu_791_p1 <= std_logic_vector(resize(unsigned(p_0554_2_fu_784_p3),3));
    p_0554_2_fu_784_p3 <= 
        sign_cnt_V_1_fu_755_p2 when (zh_2_1_V_reg_993(0) = '1') else 
        p_0554_1_fu_722_p3;
    p_0554_3_fu_801_p3 <= 
        sign_cnt_V_2_fu_795_p2 when (zh_2_2_V_reg_1002(0) = '1') else 
        p_0554_2_cast_fu_791_p1;
    p_1_17_fu_673_p3 <= 
        z1_2_V_fu_667_p2 when (tmp_36_fu_648_p1(0) = '1') else 
        z1_2_V_cast_fu_610_p1;
    p_5_cast_fu_657_p1 <= std_logic_vector(resize(unsigned(not_tmp_s_fu_652_p2),2));
    p_neg1_fu_581_p2 <= std_logic_vector(unsigned(p_neg_fu_575_p2) - unsigned(tmp_39_fu_571_p1));
    p_neg_fu_575_p2 <= std_logic_vector(unsigned(p_0622_1_reg_264) + unsigned(ap_const_lv7_70));
    p_s_16_fu_620_p3 <= 
        z1_1_V_fu_614_p2 when (tmp_35_reg_1025(0) = '1') else 
        z1_1_V_cast_fu_600_p1;
    
    zh_2_1_V_reg_993_temp <= signed(zh_2_1_V_reg_993);
    phitmp1761_s_fu_733_p1 <= std_logic_vector(resize(zh_2_1_V_reg_993_temp,2));

    phitmp1761_s_fu_733_p3 <= 
        phitmp1761_s_fu_733_p1 when (tmp_37_fu_718_p1(0) = '1') else 
        zh_2_1_V_cast_fu_587_p1;
    
    zh_2_2_V_reg_1002_temp <= signed(zh_2_2_V_reg_1002);
    phitmp1763_s_fu_818_p1 <= std_logic_vector(resize(zh_2_2_V_reg_1002_temp,2));

    phitmp1763_s_fu_818_p3 <= 
        phitmp1763_s_fu_818_p1 when (tmp_38_reg_1053(0) = '1') else 
        zh_2_2_V_cast_fu_808_p1;
    phitmp_fu_590_p4 <= lhs_V_reg_253(15 downto 8);
    r_V_10_fu_347_p2 <= (r_V_9_fu_341_p2 or lhs_V_reg_253);
    r_V_11_fu_627_p1 <= std_logic_vector(resize(unsigned(r_V_s_reg_1038),32));
    r_V_12_fu_691_p1 <= std_logic_vector(resize(unsigned(r_V_1_fu_681_p4),32));
    r_V_13_fu_751_p1 <= std_logic_vector(resize(unsigned(r_V_2_fu_741_p4),32));
    r_V_14_fu_895_p3 <= 
        tmp_28_fu_889_p2 when (tmp_40_fu_857_p3(0) = '1') else 
        tmp_25_fu_869_p2;
    r_V_1_fu_681_p4 <= signs_V_2_fu_642_p3(31 downto 1);
    r_V_2_fu_741_p4 <= signs_V_4_fu_710_p3(31 downto 1);
    r_V_9_fu_341_p2 <= std_logic_vector(shift_left(unsigned(temp_V_fu_333_p1),to_integer(unsigned('0' & tmp_7_fu_337_p1(31-1 downto 0)))));
    r_V_fu_539_p3 <= 
        tmp_20_fu_533_p2 when (tmp_33_fu_501_p3(0) = '1') else 
        tmp_17_fu_513_p2;
    sign_cnt_V_1_fu_755_p2 <= std_logic_vector(unsigned(p_0554_1_fu_722_p3) + unsigned(ap_const_lv2_1));
    sign_cnt_V_2_fu_795_p2 <= std_logic_vector(unsigned(p_0554_2_cast_fu_791_p1) + unsigned(ap_const_lv3_1));
    sign_cnt_V_fu_695_p3 <= 
        ap_const_lv2_1 when (tmp_21_reg_1030(0) = '1') else 
        ap_const_lv2_2;
    signs_V_2_fu_642_p3 <= 
        signs_V_reg_1020 when (tmp_21_reg_1030(0) = '1') else 
        r_V_11_fu_627_p1;
    signs_V_4_fu_710_p3 <= 
        signs_V_2_fu_642_p3 when (tmp_22_fu_661_p2(0) = '1') else 
        r_V_12_fu_691_p1;
    signs_V_6_fu_773_p3 <= 
        r_V_13_fu_751_p1 when (zh_2_1_V_reg_993(0) = '1') else 
        signs_V_4_fu_710_p3;
    signs_V_fu_547_p1 <= r_V_fu_539_p3(32 - 1 downto 0);
    temp_V_fu_333_p1 <= std_logic_vector(resize(unsigned(code_V_V_dout),96));
    
    inner_cnt_3_phi_fu_301_p4_temp <= signed(inner_cnt_3_phi_fu_301_p4);
    tmp_10_fu_435_p1 <= std_logic_vector(resize(inner_cnt_3_phi_fu_301_p4_temp,64));

    tmp_11_cast_fu_411_p2 <= std_logic_vector(unsigned(tmp_16_fu_407_p1) + unsigned(ap_const_lv19_7FFFF));
    tmp_11_fu_443_p4 <= val_table_q0(5 downto 4);
    tmp_13_fu_479_p3 <= (tmp_11_fu_443_p4 & tmp_32_fu_475_p1);
    tmp_14_fu_603_p3 <= (tmp_12_reg_988 & phitmp_fu_590_p4);
    
    op2_assign_fu_491_p2_temp <= signed(op2_assign_fu_491_p2);
    tmp_15_fu_509_p0 <= std_logic_vector(resize(op2_assign_fu_491_p2_temp,64));

    tmp_15_fu_509_p1 <= std_logic_vector(resize(unsigned(tmp_15_fu_509_p0),96));
    tmp_16_fu_407_p1 <= tmp_9_fu_401_p2(19 - 1 downto 0);
    tmp_17_fu_513_p2 <= std_logic_vector(shift_right(unsigned(lhs_V_reg_253),to_integer(unsigned('0' & tmp_15_fu_509_p1(31-1 downto 0)))));
    tmp_18_fu_519_p1 <= tmp_23_cast_fu_487_p1;
    tmp_18_fu_519_p2 <= std_logic_vector(unsigned(ap_const_lv10_3F0) - unsigned(tmp_18_fu_519_p1));
    
    tmp_18_fu_519_p2_temp <= signed(tmp_18_fu_519_p2);
    tmp_19_fu_529_p0 <= std_logic_vector(resize(tmp_18_fu_519_p2_temp,64));

    tmp_19_fu_529_p1 <= std_logic_vector(resize(unsigned(tmp_19_fu_529_p0),96));
    tmp_1_fu_327_p2 <= "1" when (unsigned(p_0622_1_reg_264) < unsigned(ap_const_lv7_41)) else "0";
    tmp_20_fu_533_p2 <= std_logic_vector(shift_left(unsigned(lhs_V_reg_253),to_integer(unsigned('0' & tmp_19_fu_529_p1(31-1 downto 0)))));
    tmp_21_fu_555_p2 <= "1" when (tmp_13_fu_479_p3 = ap_const_lv10_0) else "0";
    tmp_22_fu_661_p2 <= "1" when (tmp_14_fu_603_p3 = ap_const_lv10_0) else "0";
    
    e_length_V_1_fu_130_temp <= signed(e_length_V_1_fu_130);
    tmp_23_cast_fu_487_p1 <= std_logic_vector(resize(e_length_V_1_fu_130_temp,10));

    tmp_23_fu_837_p1 <= std_logic_vector(resize(unsigned(p_0554_3_reg_1058),7));
    
    op2_assign_1_fu_848_p2_temp <= signed(op2_assign_1_fu_848_p2);
    tmp_24_fu_865_p0 <= std_logic_vector(resize(op2_assign_1_fu_848_p2_temp,64));

    tmp_24_fu_865_p1 <= std_logic_vector(resize(unsigned(tmp_24_fu_865_p0),96));
    tmp_25_fu_869_p2 <= std_logic_vector(shift_right(unsigned(lhs_V_reg_253),to_integer(unsigned('0' & tmp_24_fu_865_p1(31-1 downto 0)))));
    tmp_26_fu_875_p2 <= std_logic_vector(unsigned(ap_const_lv10_0) - unsigned(op2_assign_1_fu_848_p2));
    
    tmp_26_fu_875_p2_temp <= signed(tmp_26_fu_875_p2);
    tmp_27_fu_885_p0 <= std_logic_vector(resize(tmp_26_fu_875_p2_temp,64));

    tmp_27_fu_885_p1 <= std_logic_vector(resize(unsigned(tmp_27_fu_885_p0),96));
    tmp_28_fu_889_p2 <= std_logic_vector(shift_left(unsigned(lhs_V_reg_253),to_integer(unsigned('0' & tmp_27_fu_885_p1(31-1 downto 0)))));
    tmp_2_nbreadreq_fu_134_p3 <= (0=>code_V_V_empty_n, others=>'-');
    tmp_32_fu_475_p1 <= lhs_V_reg_253(8 - 1 downto 0);
    tmp_33_fu_501_p3 <= op2_assign_fu_491_p2(9 downto 9);
    tmp_35_fu_551_p1 <= r_V_fu_539_p3(1 - 1 downto 0);
    tmp_36_fu_648_p1 <= signs_V_2_fu_642_p3(1 - 1 downto 0);
    tmp_37_fu_718_p1 <= signs_V_4_fu_710_p3(1 - 1 downto 0);
    tmp_38_fu_780_p1 <= signs_V_6_fu_773_p3(1 - 1 downto 0);
    tmp_39_fu_571_p1 <= e_length_V_1_fu_130(7 - 1 downto 0);
    tmp_3_fu_417_p2 <= (tmp_11_cast_fu_411_p2 and full_e_V_reg_934);
    tmp_40_fu_857_p3 <= op2_assign_1_fu_848_p2(9 downto 9);
    tmp_44_cast_fu_845_p1 <= std_logic_vector(resize(unsigned(p_0554_3_reg_1058),10));
    tmp_4_fu_373_p3 <= inner_cnt_2_reg_275(6 downto 6);
    tmp_5_fu_387_p1 <= std_logic_vector(resize(unsigned(inner_cnt_2_reg_275),64));
    tmp_6_fu_393_p1 <= std_logic_vector(resize(unsigned(val_table_q0),64));
    tmp_7_fu_337_p1 <= std_logic_vector(resize(unsigned(p_0622_1_reg_264),96));
    tmp_8_fu_398_p1 <= std_logic_vector(resize(unsigned(bt_cnt_V_reg_974),32));
    tmp_9_fu_401_p2 <= std_logic_vector(shift_left(unsigned(ap_const_lv32_1),to_integer(unsigned('0' & tmp_8_fu_398_p1(31-1 downto 0)))));
    tmp_V_1_fu_630_p3 <= 
        ap_const_lv11_0 when (tmp_21_reg_1030(0) = '1') else 
        p_s_16_fu_620_p3;
    tmp_V_2_fu_702_p3 <= 
        ap_const_lv11_0 when (tmp_22_fu_661_p2(0) = '1') else 
        p_1_17_fu_673_p3;
    tmp_V_3_fu_761_p3 <= 
        phitmp1761_s_fu_733_p3 when (zh_2_1_V_reg_993(0) = '1') else 
        ap_const_lv2_0;
    
    tmp_V_3_fu_761_p3_temp <= signed(tmp_V_3_fu_761_p3);
    tmp_V_4_fu_768_p1 <= std_logic_vector(resize(tmp_V_3_fu_761_p3_temp,3));

    
    tmp_V_6_fu_825_p3_temp <= signed(tmp_V_6_fu_825_p3);
    tmp_V_5_fu_832_p1 <= std_logic_vector(resize(tmp_V_6_fu_825_p3_temp,3));

    
    tmp_V_1_fu_630_p3_temp <= signed(tmp_V_1_fu_630_p3);
    tmp_V_6_cast_fu_637_p1 <= std_logic_vector(resize(tmp_V_1_fu_630_p3_temp,14));

    tmp_V_6_fu_825_p3 <= 
        phitmp1763_s_fu_818_p3 when (zh_2_2_V_reg_1002(0) = '1') else 
        ap_const_lv2_0;
    
    tmp_V_2_reg_1048_temp <= signed(tmp_V_2_reg_1048);
    tmp_V_7_cast_fu_811_p1 <= std_logic_vector(resize(tmp_V_2_reg_1048_temp,14));

    tmp_fu_321_p2 <= std_logic_vector(unsigned(cnt_reg_230) + unsigned(ap_const_lv9_1));
    tmp_s_fu_422_p2 <= "1" when (tmp_3_fu_417_p2 = dec_e_table_load_reg_969) else "0";

    -- val_table_address0 assign process. --
    val_table_address0_assign_proc : process(ap_CS_fsm, tmp_5_fu_387_p1, tmp_10_fu_435_p1)
    begin
        if ((ap_ST_st7_fsm_6 = ap_CS_fsm)) then 
            val_table_address0 <= tmp_10_fu_435_p1(6 - 1 downto 0);
        elsif ((ap_ST_st4_fsm_3 = ap_CS_fsm)) then 
            val_table_address0 <= tmp_5_fu_387_p1(6 - 1 downto 0);
        else 
            val_table_address0 <= "XXXXXX";
        end if; 
    end process;


    -- val_table_ce0 assign process. --
    val_table_ce0_assign_proc : process(ap_CS_fsm)
    begin
        if (((ap_ST_st4_fsm_3 = ap_CS_fsm) or (ap_ST_st7_fsm_6 = ap_CS_fsm))) then 
            val_table_ce0 <= ap_const_logic_1;
        else 
            val_table_ce0 <= ap_const_logic_0;
        end if; 
    end process;

    z1_1_V_cast_fu_600_p1 <= std_logic_vector(resize(unsigned(tmp_13_reg_1010),11));
    z1_1_V_fu_614_p2 <= std_logic_vector(unsigned(ap_const_lv11_0) - unsigned(z1_1_V_cast_fu_600_p1));
    z1_2_V_cast_fu_610_p1 <= std_logic_vector(resize(unsigned(tmp_14_fu_603_p3),11));
    z1_2_V_fu_667_p2 <= std_logic_vector(unsigned(ap_const_lv11_0) - unsigned(z1_2_V_cast_fu_610_p1));

    -- z1_V_V_din assign process. --
    z1_V_V_din_assign_proc : process(ap_CS_fsm, ap_sig_bdd_142, tmp_V_6_cast_fu_637_p1, tmp_V_7_cast_fu_811_p1)
    begin
        if (not(ap_sig_bdd_142)) then
            if ((ap_ST_st10_fsm_9 = ap_CS_fsm)) then 
                z1_V_V_din <= tmp_V_7_cast_fu_811_p1;
            elsif ((ap_ST_st9_fsm_8 = ap_CS_fsm)) then 
                z1_V_V_din <= tmp_V_6_cast_fu_637_p1;
            else 
                z1_V_V_din <= "XXXXXXXXXXXXXX";
            end if;
        else 
            z1_V_V_din <= "XXXXXXXXXXXXXX";
        end if; 
    end process;


    -- z1_V_V_write assign process. --
    z1_V_V_write_assign_proc : process(ap_CS_fsm, ap_sig_bdd_142)
    begin
        if ((((ap_ST_st9_fsm_8 = ap_CS_fsm) and not(ap_sig_bdd_142)) or (not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm)))) then 
            z1_V_V_write <= ap_const_logic_1;
        else 
            z1_V_V_write <= ap_const_logic_0;
        end if; 
    end process;


    -- z2_V_V_din assign process. --
    z2_V_V_din_assign_proc : process(ap_CS_fsm, ap_sig_bdd_142, tmp_V_4_fu_768_p1, tmp_V_5_fu_832_p1)
    begin
        if (not(ap_sig_bdd_142)) then
            if ((ap_ST_st10_fsm_9 = ap_CS_fsm)) then 
                z2_V_V_din <= tmp_V_5_fu_832_p1;
            elsif ((ap_ST_st9_fsm_8 = ap_CS_fsm)) then 
                z2_V_V_din <= tmp_V_4_fu_768_p1;
            else 
                z2_V_V_din <= "XXX";
            end if;
        else 
            z2_V_V_din <= "XXX";
        end if; 
    end process;


    -- z2_V_V_write assign process. --
    z2_V_V_write_assign_proc : process(ap_CS_fsm, ap_sig_bdd_142)
    begin
        if ((((ap_ST_st9_fsm_8 = ap_CS_fsm) and not(ap_sig_bdd_142)) or (not(ap_sig_bdd_142) and (ap_ST_st10_fsm_9 = ap_CS_fsm)))) then 
            z2_V_V_write <= ap_const_logic_1;
        else 
            z2_V_V_write <= ap_const_logic_0;
        end if; 
    end process;

    zh_2_1_V_cast_fu_587_p1 <= std_logic_vector(resize(unsigned(zh_2_1_V_reg_993),2));
    zh_2_2_V_cast_fu_808_p1 <= std_logic_vector(resize(unsigned(zh_2_2_V_reg_1002),2));
    zh_2_2_V_fu_471_p1 <= val_table_q0(1 - 1 downto 0);
end behav;
