--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/
-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC
-- Version: 2013.4
-- Copyright (C) 2013 Xilinx Inc. All rights reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fft_mar_12289 is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    w_in_V : IN STD_LOGIC_VECTOR (13 downto 0);
    a_in_V : IN STD_LOGIC_VECTOR (13 downto 0);
    b_in_V : IN STD_LOGIC_VECTOR (13 downto 0);
    x_add_out_V : OUT STD_LOGIC_VECTOR (13 downto 0);
    x_sub_out_V : OUT STD_LOGIC_VECTOR (13 downto 0) );
end;


architecture behav of fft_mar_12289 is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "fft_mar_12289,hls_ip_2013_4,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020clg484-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=pipeline,HLS_SYN_CLOCK=8.620000,HLS_SYN_LAT=6,HLS_SYN_TPT=1,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=0,HLS_SYN_LUT=0}";
    constant ap_true : BOOLEAN := true;
    constant ap_const_lv14_0 : STD_LOGIC_VECTOR (13 downto 0) := "00000000000000";
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv2_0 : STD_LOGIC_VECTOR (1 downto 0) := "00";
    constant ap_const_lv5_0 : STD_LOGIC_VECTOR (4 downto 0) := "00000";
    constant ap_const_lv7_0 : STD_LOGIC_VECTOR (6 downto 0) := "0000000";
    constant ap_const_lv9_0 : STD_LOGIC_VECTOR (8 downto 0) := "000000000";
    constant ap_const_lv11_0 : STD_LOGIC_VECTOR (10 downto 0) := "00000000000";
    constant ap_const_lv13_0 : STD_LOGIC_VECTOR (12 downto 0) := "0000000000000";
    constant ap_const_lv15_0 : STD_LOGIC_VECTOR (14 downto 0) := "000000000000000";
    constant ap_const_lv32_1D : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011101";
    constant ap_const_lv32_2B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101011";
    constant ap_const_lv12_0 : STD_LOGIC_VECTOR (11 downto 0) := "000000000000";
    constant ap_const_lv28_3000 : STD_LOGIC_VECTOR (27 downto 0) := "0000000000000011000000000000";
    constant ap_const_lv28_FFF : STD_LOGIC_VECTOR (27 downto 0) := "0000000000000000111111111111";
    constant ap_const_lv15_3000 : STD_LOGIC_VECTOR (14 downto 0) := "011000000000000";
    constant ap_const_lv16_FFF : STD_LOGIC_VECTOR (15 downto 0) := "0000111111111111";
    constant ap_const_lv15_3001 : STD_LOGIC_VECTOR (14 downto 0) := "011000000000001";
    constant ap_const_lv16_3000 : STD_LOGIC_VECTOR (15 downto 0) := "0011000000000000";
    constant ap_const_lv15_FFF : STD_LOGIC_VECTOR (14 downto 0) := "000111111111111";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';

    signal a_in_V_read_reg_451 : STD_LOGIC_VECTOR (13 downto 0);
    signal ap_reg_ppstg_a_in_V_read_reg_451_pp0_it1 : STD_LOGIC_VECTOR (13 downto 0);
    signal ap_reg_ppstg_a_in_V_read_reg_451_pp0_it2 : STD_LOGIC_VECTOR (13 downto 0);
    signal ap_reg_ppstg_a_in_V_read_reg_451_pp0_it3 : STD_LOGIC_VECTOR (13 downto 0);
    signal ap_reg_ppstg_a_in_V_read_reg_451_pp0_it4 : STD_LOGIC_VECTOR (13 downto 0);
    signal ap_reg_ppstg_a_in_V_read_reg_451_pp0_it5 : STD_LOGIC_VECTOR (13 downto 0);
    signal res_V_fu_135_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal res_V_reg_457 : STD_LOGIC_VECTOR (27 downto 0);
    signal ap_reg_ppstg_res_V_reg_457_pp0_it1 : STD_LOGIC_VECTOR (27 downto 0);
    signal ap_reg_ppstg_res_V_reg_457_pp0_it2 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_5_fu_184_p2 : STD_LOGIC_VECTOR (33 downto 0);
    signal r_V_5_reg_470 : STD_LOGIC_VECTOR (33 downto 0);
    signal r_V_11_fu_246_p2 : STD_LOGIC_VECTOR (39 downto 0);
    signal r_V_11_reg_475 : STD_LOGIC_VECTOR (39 downto 0);
    signal tmp_4_fu_293_p4 : STD_LOGIC_VECTOR (14 downto 0);
    signal tmp_4_reg_480 : STD_LOGIC_VECTOR (14 downto 0);
    signal p_neg_i_fu_307_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal p_neg_i_reg_486 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_7_i_fu_335_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_7_i_reg_491 : STD_LOGIC_VECTOR (27 downto 0);
    signal res_red_V_fu_358_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal res_red_V_reg_498 : STD_LOGIC_VECTOR (13 downto 0);
    signal tmp_5_fu_441_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal x_add_out_V_preg : STD_LOGIC_VECTOR (13 downto 0) := "00000000000000";
    signal tmp_8_fu_446_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal x_sub_out_V_preg : STD_LOGIC_VECTOR (13 downto 0) := "00000000000000";
    signal res_V_fu_135_p0 : STD_LOGIC_VECTOR (13 downto 0);
    signal res_V_fu_135_p1 : STD_LOGIC_VECTOR (13 downto 0);
    signal r_V_1_fu_141_p3 : STD_LOGIC_VECTOR (28 downto 0);
    signal r_V_2_fu_148_p3 : STD_LOGIC_VECTOR (29 downto 0);
    signal lhs_V_1_cast_fu_155_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal rhs_V_1_cast_fu_159_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal r_V_3_fu_163_p2 : STD_LOGIC_VECTOR (30 downto 0);
    signal r_V_4_fu_169_p3 : STD_LOGIC_VECTOR (32 downto 0);
    signal lhs_V_2_cast_fu_176_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal rhs_V_2_cast_fu_180_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal r_V_6_fu_190_p3 : STD_LOGIC_VECTOR (34 downto 0);
    signal lhs_V_3_cast_fu_197_p1 : STD_LOGIC_VECTOR (35 downto 0);
    signal rhs_V_3_cast_fu_200_p1 : STD_LOGIC_VECTOR (35 downto 0);
    signal r_V_7_fu_204_p2 : STD_LOGIC_VECTOR (35 downto 0);
    signal r_V_8_fu_210_p3 : STD_LOGIC_VECTOR (36 downto 0);
    signal lhs_V_4_cast_fu_217_p1 : STD_LOGIC_VECTOR (37 downto 0);
    signal rhs_V_4_cast_fu_221_p1 : STD_LOGIC_VECTOR (37 downto 0);
    signal r_V_9_fu_225_p2 : STD_LOGIC_VECTOR (37 downto 0);
    signal r_V_10_fu_231_p3 : STD_LOGIC_VECTOR (38 downto 0);
    signal lhs_V_5_cast_fu_238_p1 : STD_LOGIC_VECTOR (39 downto 0);
    signal rhs_V_5_cast_fu_242_p1 : STD_LOGIC_VECTOR (39 downto 0);
    signal r_V_12_fu_252_p3 : STD_LOGIC_VECTOR (40 downto 0);
    signal lhs_V_6_cast_fu_259_p1 : STD_LOGIC_VECTOR (41 downto 0);
    signal rhs_V_6_cast_fu_262_p1 : STD_LOGIC_VECTOR (41 downto 0);
    signal r_V_14_fu_272_p3 : STD_LOGIC_VECTOR (42 downto 0);
    signal r_V_13_fu_266_p2 : STD_LOGIC_VECTOR (41 downto 0);
    signal lhs_V_7_cast_fu_283_p1 : STD_LOGIC_VECTOR (43 downto 0);
    signal r_V_14_cast_fu_279_p1 : STD_LOGIC_VECTOR (43 downto 0);
    signal r_V_15_fu_287_p2 : STD_LOGIC_VECTOR (43 downto 0);
    signal phitmp_i_fu_303_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal phitmp1_i_fu_312_p3 : STD_LOGIC_VECTOR (26 downto 0);
    signal phitmp2_i_fu_323_p3 : STD_LOGIC_VECTOR (27 downto 0);
    signal p_neg1_i_fu_330_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal phitmp1_i_cast_fu_319_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_8_i_fu_341_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal p_i_fu_346_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_9_i_fu_351_p3 : STD_LOGIC_VECTOR (27 downto 0);
    signal lhs_V_fu_362_p1 : STD_LOGIC_VECTOR (14 downto 0);
    signal rhs_V_fu_365_p1 : STD_LOGIC_VECTOR (14 downto 0);
    signal r_V_fu_368_p2 : STD_LOGIC_VECTOR (14 downto 0);
    signal x_add_intern_V_fu_374_p1 : STD_LOGIC_VECTOR (15 downto 0);
    signal tmp_6_fu_378_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal x_add_intern_V_1_fu_384_p2 : STD_LOGIC_VECTOR (15 downto 0);
    signal tmp_9_fu_401_p2 : STD_LOGIC_VECTOR (14 downto 0);
    signal x_sub_intern_V_fu_411_p0 : STD_LOGIC_VECTOR (15 downto 0);
    signal tmp_9_fu_401_p2_temp: signed (15-1 downto 0);
    signal tmp_7_fu_398_p1 : STD_LOGIC_VECTOR (15 downto 0);
    signal x_sub_intern_V_fu_411_p2 : STD_LOGIC_VECTOR (15 downto 0);
    signal tmp_3_fu_417_p1 : STD_LOGIC_VECTOR (14 downto 0);
    signal tmp_s_fu_421_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal x_sub_intern_V_1_fu_427_p2 : STD_LOGIC_VECTOR (14 downto 0);
    signal x_add_intern_V_2_fu_390_p3 : STD_LOGIC_VECTOR (15 downto 0);
    signal x_sub_intern_V_2_fu_433_p3 : STD_LOGIC_VECTOR (14 downto 0);
    signal res_V_fu_135_p00 : STD_LOGIC_VECTOR (27 downto 0);
    signal res_V_fu_135_p10 : STD_LOGIC_VECTOR (27 downto 0);


begin




    -- x_add_out_V_preg assign process. --
    x_add_out_V_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                x_add_out_V_preg <= ap_const_lv14_0;
            else
                x_add_out_V_preg <= tmp_5_fu_441_p1;
            end if;
        end if;
    end process;


    -- x_sub_out_V_preg assign process. --
    x_sub_out_V_preg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                x_sub_out_V_preg <= ap_const_lv14_0;
            else
                x_sub_out_V_preg <= tmp_8_fu_446_p1;
            end if;
        end if;
    end process;


    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_true = ap_true)) then
                a_in_V_read_reg_451 <= a_in_V;
                ap_reg_ppstg_a_in_V_read_reg_451_pp0_it1 <= a_in_V_read_reg_451;
                ap_reg_ppstg_a_in_V_read_reg_451_pp0_it2 <= ap_reg_ppstg_a_in_V_read_reg_451_pp0_it1;
                ap_reg_ppstg_a_in_V_read_reg_451_pp0_it3 <= ap_reg_ppstg_a_in_V_read_reg_451_pp0_it2;
                ap_reg_ppstg_a_in_V_read_reg_451_pp0_it4 <= ap_reg_ppstg_a_in_V_read_reg_451_pp0_it3;
                ap_reg_ppstg_a_in_V_read_reg_451_pp0_it5 <= ap_reg_ppstg_a_in_V_read_reg_451_pp0_it4;
                ap_reg_ppstg_res_V_reg_457_pp0_it1 <= res_V_reg_457;
                ap_reg_ppstg_res_V_reg_457_pp0_it2 <= ap_reg_ppstg_res_V_reg_457_pp0_it1;
                p_neg_i_reg_486 <= p_neg_i_fu_307_p2;
                r_V_11_reg_475(1) <= r_V_11_fu_246_p2(1);
    r_V_11_reg_475(2) <= r_V_11_fu_246_p2(2);
    r_V_11_reg_475(3) <= r_V_11_fu_246_p2(3);
    r_V_11_reg_475(4) <= r_V_11_fu_246_p2(4);
    r_V_11_reg_475(5) <= r_V_11_fu_246_p2(5);
    r_V_11_reg_475(6) <= r_V_11_fu_246_p2(6);
    r_V_11_reg_475(7) <= r_V_11_fu_246_p2(7);
    r_V_11_reg_475(8) <= r_V_11_fu_246_p2(8);
    r_V_11_reg_475(9) <= r_V_11_fu_246_p2(9);
    r_V_11_reg_475(10) <= r_V_11_fu_246_p2(10);
    r_V_11_reg_475(11) <= r_V_11_fu_246_p2(11);
    r_V_11_reg_475(12) <= r_V_11_fu_246_p2(12);
    r_V_11_reg_475(13) <= r_V_11_fu_246_p2(13);
    r_V_11_reg_475(14) <= r_V_11_fu_246_p2(14);
    r_V_11_reg_475(15) <= r_V_11_fu_246_p2(15);
    r_V_11_reg_475(16) <= r_V_11_fu_246_p2(16);
    r_V_11_reg_475(17) <= r_V_11_fu_246_p2(17);
    r_V_11_reg_475(18) <= r_V_11_fu_246_p2(18);
    r_V_11_reg_475(19) <= r_V_11_fu_246_p2(19);
    r_V_11_reg_475(20) <= r_V_11_fu_246_p2(20);
    r_V_11_reg_475(21) <= r_V_11_fu_246_p2(21);
    r_V_11_reg_475(22) <= r_V_11_fu_246_p2(22);
    r_V_11_reg_475(23) <= r_V_11_fu_246_p2(23);
    r_V_11_reg_475(24) <= r_V_11_fu_246_p2(24);
    r_V_11_reg_475(25) <= r_V_11_fu_246_p2(25);
    r_V_11_reg_475(26) <= r_V_11_fu_246_p2(26);
    r_V_11_reg_475(27) <= r_V_11_fu_246_p2(27);
    r_V_11_reg_475(28) <= r_V_11_fu_246_p2(28);
    r_V_11_reg_475(29) <= r_V_11_fu_246_p2(29);
    r_V_11_reg_475(30) <= r_V_11_fu_246_p2(30);
    r_V_11_reg_475(31) <= r_V_11_fu_246_p2(31);
    r_V_11_reg_475(32) <= r_V_11_fu_246_p2(32);
    r_V_11_reg_475(33) <= r_V_11_fu_246_p2(33);
    r_V_11_reg_475(34) <= r_V_11_fu_246_p2(34);
    r_V_11_reg_475(35) <= r_V_11_fu_246_p2(35);
    r_V_11_reg_475(36) <= r_V_11_fu_246_p2(36);
    r_V_11_reg_475(37) <= r_V_11_fu_246_p2(37);
    r_V_11_reg_475(38) <= r_V_11_fu_246_p2(38);
    r_V_11_reg_475(39) <= r_V_11_fu_246_p2(39);
                r_V_5_reg_470(1) <= r_V_5_fu_184_p2(1);
    r_V_5_reg_470(2) <= r_V_5_fu_184_p2(2);
    r_V_5_reg_470(3) <= r_V_5_fu_184_p2(3);
    r_V_5_reg_470(4) <= r_V_5_fu_184_p2(4);
    r_V_5_reg_470(5) <= r_V_5_fu_184_p2(5);
    r_V_5_reg_470(6) <= r_V_5_fu_184_p2(6);
    r_V_5_reg_470(7) <= r_V_5_fu_184_p2(7);
    r_V_5_reg_470(8) <= r_V_5_fu_184_p2(8);
    r_V_5_reg_470(9) <= r_V_5_fu_184_p2(9);
    r_V_5_reg_470(10) <= r_V_5_fu_184_p2(10);
    r_V_5_reg_470(11) <= r_V_5_fu_184_p2(11);
    r_V_5_reg_470(12) <= r_V_5_fu_184_p2(12);
    r_V_5_reg_470(13) <= r_V_5_fu_184_p2(13);
    r_V_5_reg_470(14) <= r_V_5_fu_184_p2(14);
    r_V_5_reg_470(15) <= r_V_5_fu_184_p2(15);
    r_V_5_reg_470(16) <= r_V_5_fu_184_p2(16);
    r_V_5_reg_470(17) <= r_V_5_fu_184_p2(17);
    r_V_5_reg_470(18) <= r_V_5_fu_184_p2(18);
    r_V_5_reg_470(19) <= r_V_5_fu_184_p2(19);
    r_V_5_reg_470(20) <= r_V_5_fu_184_p2(20);
    r_V_5_reg_470(21) <= r_V_5_fu_184_p2(21);
    r_V_5_reg_470(22) <= r_V_5_fu_184_p2(22);
    r_V_5_reg_470(23) <= r_V_5_fu_184_p2(23);
    r_V_5_reg_470(24) <= r_V_5_fu_184_p2(24);
    r_V_5_reg_470(25) <= r_V_5_fu_184_p2(25);
    r_V_5_reg_470(26) <= r_V_5_fu_184_p2(26);
    r_V_5_reg_470(27) <= r_V_5_fu_184_p2(27);
    r_V_5_reg_470(28) <= r_V_5_fu_184_p2(28);
    r_V_5_reg_470(29) <= r_V_5_fu_184_p2(29);
    r_V_5_reg_470(30) <= r_V_5_fu_184_p2(30);
    r_V_5_reg_470(31) <= r_V_5_fu_184_p2(31);
    r_V_5_reg_470(32) <= r_V_5_fu_184_p2(32);
    r_V_5_reg_470(33) <= r_V_5_fu_184_p2(33);
                res_V_reg_457 <= res_V_fu_135_p2;
                res_red_V_reg_498 <= res_red_V_fu_358_p1;
                tmp_4_reg_480 <= r_V_15_fu_287_p2(43 downto 29);
                tmp_7_i_reg_491 <= tmp_7_i_fu_335_p2;
            end if;
        end if;
    end process;
    r_V_5_reg_470(0) <= '0';
    r_V_11_reg_475(0) <= '0';
    lhs_V_1_cast_fu_155_p1 <= std_logic_vector(resize(unsigned(r_V_1_fu_141_p3),31));
    lhs_V_2_cast_fu_176_p1 <= std_logic_vector(resize(unsigned(r_V_3_fu_163_p2),34));
    lhs_V_3_cast_fu_197_p1 <= std_logic_vector(resize(unsigned(r_V_5_reg_470),36));
    lhs_V_4_cast_fu_217_p1 <= std_logic_vector(resize(unsigned(r_V_7_fu_204_p2),38));
    lhs_V_5_cast_fu_238_p1 <= std_logic_vector(resize(unsigned(r_V_9_fu_225_p2),40));
    lhs_V_6_cast_fu_259_p1 <= std_logic_vector(resize(unsigned(r_V_11_reg_475),42));
    lhs_V_7_cast_fu_283_p1 <= std_logic_vector(resize(unsigned(r_V_13_fu_266_p2),44));
    lhs_V_fu_362_p1 <= std_logic_vector(resize(unsigned(ap_reg_ppstg_a_in_V_read_reg_451_pp0_it5),15));
    p_i_fu_346_p2 <= std_logic_vector(unsigned(tmp_7_i_reg_491) + unsigned(ap_const_lv28_FFF));
    p_neg1_i_fu_330_p2 <= std_logic_vector(unsigned(p_neg_i_reg_486) - unsigned(phitmp2_i_fu_323_p3));
    p_neg_i_fu_307_p2 <= std_logic_vector(unsigned(ap_reg_ppstg_res_V_reg_457_pp0_it2) - unsigned(phitmp_i_fu_303_p1));
    phitmp1_i_cast_fu_319_p1 <= std_logic_vector(resize(unsigned(phitmp1_i_fu_312_p3),28));
    phitmp1_i_fu_312_p3 <= (tmp_4_reg_480 & ap_const_lv12_0);
    phitmp2_i_fu_323_p3 <= (tmp_4_reg_480 & ap_const_lv13_0);
    phitmp_i_fu_303_p1 <= std_logic_vector(resize(unsigned(tmp_4_fu_293_p4),28));
    r_V_10_fu_231_p3 <= (ap_reg_ppstg_res_V_reg_457_pp0_it1 & ap_const_lv11_0);
    r_V_11_fu_246_p2 <= std_logic_vector(unsigned(lhs_V_5_cast_fu_238_p1) + unsigned(rhs_V_5_cast_fu_242_p1));
    r_V_12_fu_252_p3 <= (ap_reg_ppstg_res_V_reg_457_pp0_it2 & ap_const_lv13_0);
    r_V_13_fu_266_p2 <= std_logic_vector(unsigned(lhs_V_6_cast_fu_259_p1) + unsigned(rhs_V_6_cast_fu_262_p1));
    r_V_14_cast_fu_279_p1 <= std_logic_vector(resize(unsigned(r_V_14_fu_272_p3),44));
    r_V_14_fu_272_p3 <= (ap_reg_ppstg_res_V_reg_457_pp0_it2 & ap_const_lv15_0);
    r_V_15_fu_287_p2 <= std_logic_vector(unsigned(lhs_V_7_cast_fu_283_p1) + unsigned(r_V_14_cast_fu_279_p1));
    r_V_1_fu_141_p3 <= (res_V_reg_457 & ap_const_lv1_0);
    r_V_2_fu_148_p3 <= (res_V_reg_457 & ap_const_lv2_0);
    r_V_3_fu_163_p2 <= std_logic_vector(unsigned(lhs_V_1_cast_fu_155_p1) + unsigned(rhs_V_1_cast_fu_159_p1));
    r_V_4_fu_169_p3 <= (res_V_reg_457 & ap_const_lv5_0);
    r_V_5_fu_184_p2 <= std_logic_vector(unsigned(lhs_V_2_cast_fu_176_p1) + unsigned(rhs_V_2_cast_fu_180_p1));
    r_V_6_fu_190_p3 <= (ap_reg_ppstg_res_V_reg_457_pp0_it1 & ap_const_lv7_0);
    r_V_7_fu_204_p2 <= std_logic_vector(unsigned(lhs_V_3_cast_fu_197_p1) + unsigned(rhs_V_3_cast_fu_200_p1));
    r_V_8_fu_210_p3 <= (ap_reg_ppstg_res_V_reg_457_pp0_it1 & ap_const_lv9_0);
    r_V_9_fu_225_p2 <= std_logic_vector(unsigned(lhs_V_4_cast_fu_217_p1) + unsigned(rhs_V_4_cast_fu_221_p1));
    r_V_fu_368_p2 <= std_logic_vector(unsigned(lhs_V_fu_362_p1) + unsigned(rhs_V_fu_365_p1));
    res_V_fu_135_p0 <= res_V_fu_135_p00(14 - 1 downto 0);
    res_V_fu_135_p00 <= std_logic_vector(resize(unsigned(b_in_V),28));
    res_V_fu_135_p1 <= res_V_fu_135_p10(14 - 1 downto 0);
    res_V_fu_135_p10 <= std_logic_vector(resize(unsigned(w_in_V),28));
    res_V_fu_135_p2 <= std_logic_vector(resize(unsigned(res_V_fu_135_p0) * unsigned(res_V_fu_135_p1), 28));
    res_red_V_fu_358_p1 <= tmp_9_i_fu_351_p3(14 - 1 downto 0);
    rhs_V_1_cast_fu_159_p1 <= std_logic_vector(resize(unsigned(r_V_2_fu_148_p3),31));
    rhs_V_2_cast_fu_180_p1 <= std_logic_vector(resize(unsigned(r_V_4_fu_169_p3),34));
    rhs_V_3_cast_fu_200_p1 <= std_logic_vector(resize(unsigned(r_V_6_fu_190_p3),36));
    rhs_V_4_cast_fu_221_p1 <= std_logic_vector(resize(unsigned(r_V_8_fu_210_p3),38));
    rhs_V_5_cast_fu_242_p1 <= std_logic_vector(resize(unsigned(r_V_10_fu_231_p3),40));
    rhs_V_6_cast_fu_262_p1 <= std_logic_vector(resize(unsigned(r_V_12_fu_252_p3),42));
    rhs_V_fu_365_p1 <= std_logic_vector(resize(unsigned(res_red_V_reg_498),15));
    tmp_3_fu_417_p1 <= x_sub_intern_V_fu_411_p2(15 - 1 downto 0);
    tmp_4_fu_293_p4 <= r_V_15_fu_287_p2(43 downto 29);
    tmp_5_fu_441_p1 <= x_add_intern_V_2_fu_390_p3(14 - 1 downto 0);
    tmp_6_fu_378_p2 <= "1" when (unsigned(r_V_fu_368_p2) > unsigned(ap_const_lv15_3000)) else "0";
    tmp_7_fu_398_p1 <= std_logic_vector(resize(unsigned(ap_reg_ppstg_a_in_V_read_reg_451_pp0_it5),16));
    tmp_7_i_fu_335_p2 <= std_logic_vector(unsigned(p_neg1_i_fu_330_p2) - unsigned(phitmp1_i_cast_fu_319_p1));
    tmp_8_fu_446_p1 <= x_sub_intern_V_2_fu_433_p3(14 - 1 downto 0);
    tmp_8_i_fu_341_p2 <= "1" when (unsigned(tmp_7_i_reg_491) > unsigned(ap_const_lv28_3000)) else "0";
    tmp_9_fu_401_p2 <= std_logic_vector(unsigned(ap_const_lv15_3001) - unsigned(rhs_V_fu_365_p1));
    tmp_9_i_fu_351_p3 <= 
        p_i_fu_346_p2 when (tmp_8_i_fu_341_p2(0) = '1') else 
        tmp_7_i_reg_491;
    tmp_s_fu_421_p2 <= "1" when (unsigned(x_sub_intern_V_fu_411_p2) > unsigned(ap_const_lv16_3000)) else "0";
    x_add_intern_V_1_fu_384_p2 <= std_logic_vector(unsigned(x_add_intern_V_fu_374_p1) + unsigned(ap_const_lv16_FFF));
    x_add_intern_V_2_fu_390_p3 <= 
        x_add_intern_V_1_fu_384_p2 when (tmp_6_fu_378_p2(0) = '1') else 
        x_add_intern_V_fu_374_p1;
    x_add_intern_V_fu_374_p1 <= std_logic_vector(resize(unsigned(r_V_fu_368_p2),16));

    -- x_add_out_V assign process. --
    x_add_out_V_assign_proc : process(tmp_5_fu_441_p1, x_add_out_V_preg)
    begin
        x_add_out_V <= tmp_5_fu_441_p1;
    end process;

    x_sub_intern_V_1_fu_427_p2 <= std_logic_vector(unsigned(tmp_3_fu_417_p1) + unsigned(ap_const_lv15_FFF));
    x_sub_intern_V_2_fu_433_p3 <= 
        x_sub_intern_V_1_fu_427_p2 when (tmp_s_fu_421_p2(0) = '1') else 
        tmp_3_fu_417_p1;
    
    tmp_9_fu_401_p2_temp <= signed(tmp_9_fu_401_p2);
    x_sub_intern_V_fu_411_p0 <= std_logic_vector(resize(tmp_9_fu_401_p2_temp,16));

    x_sub_intern_V_fu_411_p2 <= std_logic_vector(unsigned(x_sub_intern_V_fu_411_p0) + unsigned(tmp_7_fu_398_p1));

    -- x_sub_out_V assign process. --
    x_sub_out_V_assign_proc : process(tmp_8_fu_446_p1, x_sub_out_V_preg)
    begin
        x_sub_out_V <= tmp_8_fu_446_p1;
    end process;

end behav;
