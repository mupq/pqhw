--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:13:05 02/03/2014 
-- Design Name: 
-- Module Name:    ber_eval - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.ber_sampler_pkg.all;


--XXX TODO: Maybe split up the ROM into smaller tables. Then access should be
--cheaper and simpler. Use then a distributed RAM. This RAM can also be shared
--with other modules.
--Currently no memory LUTs are used which impacts performance and area usage


entity ber_eval is
  generic (
    PARAM_SET : integer := 1;
    MAX_PREC  : integer := 79;
    CONST_K   : integer := 253;
    MAX_X     : integer := 10
    );
  port (
    clk : in std_logic;

    rejected_value : out std_logic := '0';


    --Fifo interface to get randomness
    rand_rd_en : out std_logic;
    rand_din   : in  std_logic;
    rand_empty : in  std_logic;
    rand_valid : in  std_logic;

    fifo_ber_empty : in  std_logic;
    fifo_ber_rd_en : out std_logic;
    fifo_ber_valid : in  std_logic;
    fifo_ber_in    : in  std_logic_vector(integer(ceil(log2(real((CONST_K-1)*((CONST_K-1)+2*CONST_K*MAX_X)))))-1 downto 0);
    fifo_z_empty   : in  std_logic;
    fifo_z_rd_en   : out std_logic;
    fifo_z_valid   : in  std_logic;
    fifo_z_in      : in  std_logic_vector(integer(ceil(log2(real((CONST_K)*(MAX_X)+CONST_K-1))))-1 downto 0);

    z_dout  : out std_logic_vector(integer(ceil(log2(real((CONST_K)*(MAX_X)+CONST_K-1))))-1 downto 0) := (others => '0');
    z_full  : in  std_logic;
    z_wr_en : out std_logic
    );
end ber_eval;

architecture Behavioral of ber_eval is

  constant MAX_BER : integer := fifo_ber_in'length;
  constant MAX_Z   : integer := fifo_z_in'length;


  --constant bernoulli_vals : bernoulli_vals_type := (
  --  "1111111111111111010010100101001001111000111011101000010110111000100011100111001",
  --  "1111111111111110100101001010010101110010110010111110001000001111101010001011001",
  --  "1111111111111101001010010100110011101001010100011011000010011000101101001101010",
  --  "1111111111111010010100101010000111100001011111111010001100011110110011011100101",
  --  "1111111111110100101001010110001111111110000101001100111100010101001000111101000",
  --  "1111111111101001010010110100100011100101101000111101100011001100001100001101111",
  --  "1111111111010010100110001001010101011010010100100011100101110111011010000011110",
  --  "1111111110100101001110010011100000111001111010011010111111000110000100010110001",
  --  "1111111101001010100100101010000011010010101001000100100110001100100111111001010",
  --  "1111111010010101101001011101010101111100100110001110011011001100000010011100011",
  --  "1111110100101101010011001000111000011001001011110101100010011111001110011000001",
  --  "1111101001100010100100010101010011011110101000010001110110100011111011110100011",
  --  "1111010011100100101010011100110101011010010011100110000110010100001111111100010",
  --  "1110101001000100101011111110111001011010100011110000101110010101101001111101100",
  --  "1101011001100001101001000000110110101101000101010101101011100111110100100011010",
  --  "1011001110000111011000111000010010011000110111100110010010101000110111001100011",
  --  "0111110111100110100111001100010110001010010100000000111000111100010100010101001",
  --  "0011110111101011000001001101011011111100000010000000111011000000001101110001011",
  --  "0000111011111001110110000001000001010110111001011111101000111101010001010011010",
  --  "0000000011100000010001110111011111001111101001011100011001101110100011110100100",
  --  "0000000000000000110001000111110100100101100111110000111101011011111010100001100",
  --  "0000000000000000000000000000000010010110110011111101111011001001010100100110000");

  ----"0000000000000000000000000000000000000000000000000000000000000000010110001101100");
  type bernoulli_vals_type_80 is array (natural range <>) of std_logic_vector(128-1 downto 0);
  constant bernoulli_vals_param_1 : bernoulli_vals_type_80 := (
    "11111111111111110100101110111111111101110101111000011110001100111001001111110110010110010011101101100100000010111010111111010101",
    "11111111111111101001011110000000011011011010011001011000100011110001111010101111100101010001010011110000011110001011010011111110",
    "11111111111111010010111100000010110101101111001110111100010011001110110011101011001010000011111000110110011100010111011001111110",
    "11111111111110100101111000001101100111000111100001111001110110001111111101111000010110100000101100101000100001010010000000011000",
    "11111111111101001011110000111010111100101101101110011101101011100000011000011111100000110100101101011001101001101011100011011000",
    "11111111111010010111100011110100110010101001011100011001000010101100010101101101011100011111111110011111110011000010101111010110",
    "11111111110100101111001111100101000100100101100000110010111011111000001011000000000011001010011101000011111000110101000000011011",
    "11111111101001011110111110110111011001101011101001111011111110011111101100111011011101001000111100111100011101011011110110100000",
    "11111111010010111111111100011110010000011000100111100100100101000000111000010001011100011111101101100101001110010011011000000101",
    "11111110100110000111110011001101110000001000100001100110010011110000010100111110110101100101111101001011110100101100110011110100",
    "11111101001100101111001001111100101110110011101101000100111000000101101010011100001101011100101001010110101001101110010000000010",
    "11111010011011011011110101101110001010000111110001011000000011000101001101001110101100000101011010100101101010000100111100001100",
    "11110100111110101000010100000110000000110000110100101101000010010111100001111001100101101110111001110001100101110000101111111100",
    "11101010011011101000001010111011100010101010111001010010111001011101100110011010010110001000110100100010011110100000100110101000",
    "11010110101011100011011010110011011101010111010011011111100110000110000101010100000111110110011101011111101000111011001011001011",
    "10110100000001111011101000000010011100000000001101000100000011010111101110000101111101001011111111001011101010010010010110010001",
    "01111110100110101101110111001111001000001100111001000010101010110101111001100100101001001100110000100101000111101100110010100110",
    "00111110100111001101000000000111100000011010110111001000000000110001011111111000100011000100010111011010001100111101011101001100",
    "00001111010100000101010011010001110101010000001001101011101000000000000110011000001010111000011100001100111101111111001010100111",
    "00000000111010101000001100100101101101100011010111001001111001110001101000000010100101111010000110011101010110110100000010010011",
    "00000000000000001101011011010100000001000010000010111000010111100101010001011010111101001000101100110001010011000001001010111001",
    "00000000000000000000000000000000101101000100011100100110011111011000101010000000000110110011010101010110011111010110011101011011"
    );

  constant bernoulli_vals_param_3 : bernoulli_vals_type_80 := (
"11111111111111110111101001011111000100001000000000001110110000110011110001011010101001101011111111001101001001111010011101110011",
"11111111111111101111010010111110011001101100000010111011100011011010100101011100001000010001111010101010101001111110010101111001",
"11111111111111011110100101111101111001001000001101011101100101000111100101011100001101000111101010010101100101000111011110001110",
"11111111111110111101001100000000001001010000100111000111111101001101010111011001011110101100110110101100001100010111100111000010",
"11111111111101111010011000010001101110011111101101011010100101100000000100011100000001111100110101111101111111111011100011011010",
"11111111111011110100110001101001001100100111001010011111111010111101011110100101110011001011011001111111001100101001111101010111",
"11111111110111101001100111101001010101011011101100101101110011001110110011100101001001101011010000010111111001100100010111110110",
"11111111101111010011100000101110001001100000010001010011000010001001011110001001100010000000000100010000001111011101110011110100",
"11111111011110101000000111000111111100000011010011111000110000010100110000011010101000000010000011010001000010101011010000111101",
"11111110111101010100100100101100010001001110010110010110010010101110010001001010011111001111100110010101011100001000001101101101",
"11111101111010111010100000111000111111000101110110111100101000001111100110001001111011000100000101110010101001000111010001000111",
"11111011110110111010001101101110111010011111101101110010110110001110011000100011001110111101001011010010011010000111010111101110",
"11110111110010000110111011101100100001101110110111010101011011111111000010010101011011010001011110100011100010000000011111010011",
"11101111110101000110001011111001111011100000000111100011111110001111001000110011110100111000100000100010110101001101000111110000",
"11100000101011100100000100000010101111101001111000001001000001101011100000001101100000100110101111010110100101100111101101010000",
"11000101001100010110100001100001001111011101001000010011011100111101000000110110010110110010000011011100011000001001000001100110",
"10010111111001010001010000101110110010001110111000100011100001100100100010110111111111011010100010000101101100101010001100010011",
"01011010001000000000101011001100010011100101001110111111111001100000000011011101110110110000111101100011001101100001110000110001",
"00011111101110101000101110011010010110101001101100010001000010010010101010001011001010000111011001110011110100011111001011101010",
"00000011111011101011010110111110100010100101111000110010111010101000000011000001010111110010010111011101101100000000101100100011",
"00000000000011110111011011011000111001101000111001111001110100110000110110101000110011110111111010011110010101101001010011111001",
"00000000000000000000000011101111001001001001011110110001000000110111111100011100000100001011100110011001101001010001101011001111"
);

  constant bernoulli_vals_param_4 : bernoulli_vals_type_80 := (
"11111111111111111000111001101111011001100000001010001101010101111001011000101010000100100100011000000110110111001011101010000101",
"11111111111111110001110011011110111111100110011000010100010011101000010101001110101111010110101100011101000000000110100001000001",
"11111111111111100011100110111110110001100100111110110101101101010110110001001011100011101001000100101101111000010110001000101001",
"11111111111111000111001110000000101100101010101011010100101001100111100010011101010101010110000011010001100110100001010110011011",
"11111111111110001110011100001101111111010110110011110101001011101110111010011011000111100110001110001101101011110001101100111101",
"11111111111100011100111001001110010110101000010001010011101011001110010010110011011101110111001111101111110010001110010110011010",
"11111111111000111001110101100110001011100001110000111101100000000011101001110010101011101000100000001000000010101010110001011000",
"11111111110001110011110111110010000100111101100010000101111100011111000000010110100100100010101101011010100011011101000001101101",
"11111111100011101000100001111001101000001110000101110111110101101111000100101100100111110010001010000010001000000001100010111010",
"11111111000111010100001100111101111111100011000100011011100110000011000001111100101110000101011100111100001011001010010111001010",
"11111110001110110100111101001101110011100001101011101110001010100100010101010001101111111001010110000101000001011001100110110111",
"11111100011110011011111100011100000010110110101110001101110111111110101000101010111000100011001001110000000001100011101001110111",
"11111000111111111110101000100101011011011010100101100111000110011111000001101101010111011010010101111101000100001100001001000110",
"11110010001100001101010101111100110100010011000100100001001100000011100111101101110010100011111000000001010100011010111010000001",
"11100101001000000101110011110000101111000101100001000110001000101011001101011110111101000100010101011001111111111111000000010111",
"11001101000100101110101001011110000011101110001011101101010011001100000000010010111100000011000011111000011111000000010100011000",
"10100100010001110100110011000000011011111010000110011101101111000001001110111101100001011111010000011110010101111110001000101111",
"01101001011010110110111000110010001110001100011111010000101011100001000001011111100110010110100000011000111110101011011110101101",
"00101011011010010100110101111010011111111111111010010010110111010010110011101011001111010001010001101110100100101000011100010110",
"00000111010111001000101101010111110011001110111101101111110010000010100110000001011110100011000010000000100100111111111101001100",
"00000000001101100011000100010011010000000010100011011010110111100011110001010010101110101111011000110101010010010100010111101100",
"00000000000000000000101101111000101111011000011101110001001111101000111110101111011101101110111110111110011100111111001011011010",
"00000000000000000000000000000000000000001000001110011001001110111101111100000110110011111101111011001010111101010000010111110000"
);

  
  signal ber_val : std_logic_vector(MAX_BER-1 downto 0) := (others => '0');
  signal z_val   : std_logic_vector(MAX_Z-1 downto 0)   := (others => '0');


  signal z_val_out  : std_logic_vector(MAX_Z-1 downto 0) := (others => '0');
  signal z_val_free : std_logic                          := '1';

  signal bernoulli_line : std_logic_vector(MAX_PREC-1 downto 0) := (others => '0');
  signal counter_exp    : integer range 0 to MAX_BER-1          := 0;
  signal counter_ber    : integer range 0 to MAX_PREC-1         := 0;

  type   eg_state is (IDLE, WAIT_RAND, WAIT_RAND2, STORE, BERNOULLI, REJECTION, FIN, WAIT_RAND_AVAIL, WAIT_CYCLE);
  signal state_reg : eg_state := IDLE;

  signal read_once : std_logic := '1';

  signal bernoulli_bit     : std_logic                    := '1';
  signal bernoulli_bit_std : std_logic_vector(0 downto 0) := "0";

  signal next_one          : integer range -1 to MAX_BER-1 := 0;
  signal rand_rd_en_intern : std_logic                     := '0';

  signal sample_counter : integer := 0;

  

begin




  process (ber_val, counter_exp)
  begin  -- process
    next_one <= -1;
    for i in 0 to fifo_ber_in'length-1 loop
      if ber_val(i) = '1' and i <= counter_exp then
        next_one <= i;
      end if;
    end loop;  -- i
  end process;

  bernoulli_bit <= bernoulli_line(counter_ber);
  --bernoulli_bit_std <=std_logic_vector( resize(unsigned(bernoulli_line) srl counter_ber,1));
  --bernoulli_bit <= bernoulli_bit_std(0);

  --fifo_ber_rd_en <= '1' when (fifo_ber_empty = '0' and fifo_z_empty = '0' and state_reg = IDLE) else '0';
  --fifo_z_rd_en   <= '1' when (fifo_ber_empty = '0' and fifo_z_empty = '0' and state_reg = IDLE) else '0';

  rand_rd_en <= '1' when (state_reg = BERNOULLI and next_one /= -1 and rand_empty = '0') else rand_rd_en_intern;


  process(clk)
  begin  -- process c
    if rising_edge(clk) then
      rejected_value <= '0';

      if next_one >= 0 then
        if PARAM_SET = 1 then
          bernoulli_line <= bernoulli_vals_param_1(next_one);
        elsif PARAM_SET = 3 then
          bernoulli_line <= bernoulli_vals_param_3(next_one);
        elsif PARAM_SET = 4 then
          bernoulli_line <= bernoulli_vals_param_4(next_one);
        end if;

      end if;


      z_wr_en           <= '0';
      fifo_ber_rd_en    <= '0';
      fifo_z_rd_en      <= '0';
      rand_rd_en_intern <= '0';



      case state_reg is
        when IDLE =>
          if fifo_ber_empty = '0' and fifo_z_empty = '0' then
            fifo_ber_rd_en <= '1';
            fifo_z_rd_en   <= '1';
            state_reg      <= WAIT_CYCLE;
            --state_reg <= STORE;
          end if;

        when WAIT_CYCLE =>
          state_reg <= STORE;

          
        when STORE =>
          --Store both values in a register
          if fifo_z_valid = '1' and fifo_ber_valid = '1' then
            ber_val     <= fifo_ber_in;
            z_val       <= fifo_z_in;
            counter_exp <= MAX_BER-1;
            state_reg   <= BERNOULLI;
            z_wr_en     <= '0';
          else
            state_reg <= IDLE;
          end if;


        when BERNOULLI =>
          if rand_empty = '0' then
            if next_one = -1 then
              --If there is no more onw, then we are finished
              state_reg <= FIN;
            else
              --A one has been found
              counter_exp <= next_one;
              --state_reg         <= WAIT_RAND;
              state_reg   <= REJECTION;
              --rand_rd_en_intern <= '1';
              counter_ber <= MAX_PREC-1;
            end if;
          end if;


          --when BERNOULLI =>
          --  --Do the rejection sampling
          --  --There should be randomness available
          --  if rand_empty = '0' then
          --    --Whole poly has been checked -> Finished
          --    --See if a one bit is set, then do rejection sampling
          --    if ber_val(counter_exp) = '1' then
          --      rand_rd_en  <= '1';
          --      state_reg   <= WAIT_RAND;
          --      counter_ber <= MAX_PREC-1;
          --    else
          --      --Some more logic, to search for zer
          --      if counter_exp > 2 then
          --        if ber_val(counter_exp-1) = '0' then
          --          counter_exp <= counter_exp-2;
          --        else
          --          counter_exp <= counter_exp-1;
          --          rand_rd_en  <= '1';
          --          state_reg   <= WAIT_RAND;
          --          counter_ber <= MAX_PREC-1;
          --        end if;
          --      else
          --        if counter_exp > 0 then
          --          counter_exp <= counter_exp-1;
          --        elsif counter_exp = 0 then
          --          --The last bit is not one, we can accept
          --          state_reg <= FIN;
          --        end if;
          --      end if;
          --    end if;
          --  end if;


        when WAIT_RAND =>
          state_reg <= REJECTION;

        when REJECTION =>
          if rand_valid = '1' then
            if (bernoulli_bit = '1' and rand_din = '1') or (bernoulli_bit = '0' and rand_din = '0') then
              --Nothing happened - no decision made
              counter_ber <= counter_ber-1;

              if rand_empty = '1' then
                state_reg <= WAIT_RAND_AVAIL;
              else
                state_reg         <= WAIT_RAND2;
                rand_rd_en_intern <= '1';
              end if;

            elsif bernoulli_bit = '1' and rand_din = '0' then
              --smaller = accept this line. See next lines
              state_reg <= BERNOULLI;
              if counter_exp = 0 then
                state_reg <= FIN;
              else
                counter_exp <= counter_exp-1;
              end if;
            elsif bernoulli_bit = '0' and rand_din = '1' then
              --greater = reject
              rejected_value <= '1';
              state_reg      <= IDLE;
            end if;
          end if;

        when WAIT_RAND_AVAIL =>
          if rand_empty = '0' then
            state_reg         <= WAIT_RAND2;
            rand_rd_en_intern <= '1';
          end if;

        when WAIT_RAND2 =>
          state_reg <= REJECTION;

        when FIN =>
          --Final buffer
          -- if z_full = '0' and z_val_free = '0' then
          --   z_dout         <= z_val_out;
          --   z_wr_en        <= '1';
          --   z_val_free     <= '1';
          --   sample_counter <= sample_counter+1;
          -- end if;

          if z_full = '0' then
            state_reg <= IDLE;
            z_dout    <= z_val;
            z_wr_en   <= '1';
          end if;

          
      end case;
    end if;
  end process;


end Behavioral;





----constant bernoulli_vals : bernoulli_vals_type := (
----  "1111111111111111010010100101001001111000111011101000010110111000100011100111001",
----  "1111111111111110100101001010010101110010110010111110001000001111101010001011001",
----  "1111111111111101001010010100110011101001010100011011000010011000101101001101010",
----  "1111111111111010010100101010000111100001011111111010001100011110110011011100101",
----  "1111111111110100101001010110001111111110000101001100111100010101001000111101000",
----  "1111111111101001010010110100100011100101101000111101100011001100001100001101111",
----  "1111111111010010100110001001010101011010010100100011100101110111011010000011110",
----  "1111111110100101001110010011100000111001111010011010111111000110000100010110001",
----  "1111111101001010100100101010000011010010101001000100100110001100100111111001010",
----  "1111111010010101101001011101010101111100100110001110011011001100000010011100011",
----  "1111110100101101010011001000111000011001001011110101100010011111001110011000001",
----  "1111101001100010100100010101010011011110101000010001110110100011111011110100011",
----  "1111010011100100101010011100110101011010010011100110000110010100001111111100010",
----  "1110101001000100101011111110111001011010100011110000101110010101101001111101100",
----  "1101011001100001101001000000110110101101000101010101101011100111110100100011010",
----  "1011001110000111011000111000010010011000110111100110010010101000110111001100011",
----  "0111110111100110100111001100010110001010010100000000111000111100010100010101001",
----  "0011110111101011000001001101011011111100000010000000111011000000001101110001011",
----  "0000111011111001110110000001000001010110111001011111101000111101010001010011010",
----  "0000000011100000010001110111011111001111101001011100011001101110100011110100100",
----  "0000000000000000110001000111110100100101100111110000111101011011111010100001100",
----  "0000000000000000000000000000000010010110110011111101111011001001010100100110000");

------"0000000000000000000000000000000000000000000000000000000000000000010110001101100");
--type bernoulli_vals_type_80 is array (natural range <>) of std_logic_vector(80-1 downto 0);
--constant bernoulli_vals_param_1 : bernoulli_vals_type_80 := (
--  "11111111111111110100101110111111111101110101111000011110001100111001001111110110",
--  "11111111111111101001011110000000011011011010011001011000100011110001111010101111",
--  "11111111111111010010111100000010110101101111001110111100010011001110110011101011",
--  "11111111111110100101111000001101100111000111100001111001110110001111111101111000",
--  "11111111111101001011110000111010111100101101101110011101101011100000011000011111",
--  "11111111111010010111100011110100110010101001011100011001000010101100010101101101",
--  "11111111110100101111001111100101000100100101100000110010111011111000001011000000",
--  "11111111101001011110111110110111011001101011101001111011111110011111101100111011",
--  "11111111010010111111111100011110010000011000100111100100100101000000111000010001",
--  "11111110100110000111110011001101110000001000100001100110010011110000010100111110",
--  "11111101001100101111001001111100101110110011101101000100111000000101101010011100",
--  "11111010011011011011110101101110001010000111110001011000000011000101001101001110",
--  "11110100111110101000010100000110000000110000110100101101000010010111100001111001",
--  "11101010011011101000001010111011100010101010111001010010111001011101100110011010",
--  "11010110101011100011011010110011011101010111010011011111100110000110000101010100",
--  "10110100000001111011101000000010011100000000001101000100000011010111101110000101",
--  "01111110100110101101110111001111001000001100111001000010101010110101111001100100",
--  "00111110100111001101000000000111100000011010110111001000000000110001011111111000",
--  "00001111010100000101010011010001110101010000001001101011101000000000000110011000",
--  "00000000111010101000001100100101101101100011010111001001111001110001101000000010",
--  "00000000000000001101011011010100000001000010000010111000010111100101010001011010",
--  "00000000000000000000000000000000101101000100011100100110011111011000101010000000");

--constant bernoulli_vals_param_3 : bernoulli_vals_type_80 := (
--  "11111111111111110111101001011111000100001000000000001110110000110011110001011010",
--  "11111111111111101111010010111110011001101100000010111011100011011010100101011100",
--  "11111111111111011110100101111101111001001000001101011101100101000111100101011100",
--  "11111111111110111101001100000000001001010000100111000111111101001101010111011001",
--  "11111111111101111010011000010001101110011111101101011010100101100000000100011100",
--  "11111111111011110100110001101001001100100111001010011111111010111101011110100101",
--  "11111111110111101001100111101001010101011011101100101101110011001110110011100101",
--  "11111111101111010011100000101110001001100000010001010011000010001001011110001001",
--  "11111111011110101000000111000111111100000011010011111000110000010100110000011010",
--  "11111110111101010100100100101100010001001110010110010110010010101110010001001010",
--  "11111101111010111010100000111000111111000101110110111100101000001111100110001001",
--  "11111011110110111010001101101110111010011111101101110010110110001110011000100011",
--  "11110111110010000110111011101100100001101110110111010101011011111111000010010101",
--  "11101111110101000110001011111001111011100000000111100011111110001111001000110011",
--  "11100000101011100100000100000010101111101001111000001001000001101011100000001101",
--  "11000101001100010110100001100001001111011101001000010011011100111101000000110110",
--  "10010111111001010001010000101110110010001110111000100011100001100100100010110111",
--  "01011010001000000000101011001100010011100101001110111111111001100000000011011101",
--  "00011111101110101000101110011010010110101001101100010001000010010010101010001011",
--  "00000011111011101011010110111110100010100101111000110010111010101000000011000001",
--  "00000000000011110111011011011000111001101000111001111001110100110000110110101000",
--  "00000000000000000000000011101111001001001001011110110001000000110111111100011100");

--constant bernoulli_vals_param_4 : bernoulli_vals_type_80 := (
--  "11111111111111111000111001101111011001100000001010001101010101111001011000101010",
--  "11111111111111110001110011011110111111100110011000010100010011101000010101001110",
--  "11111111111111100011100110111110110001100100111110110101101101010110110001001011",
--  "11111111111111000111001110000000101100101010101011010100101001100111100010011101",
--  "11111111111110001110011100001101111111010110110011110101001011101110111010011011",
--  "11111111111100011100111001001110010110101000010001010011101011001110010010110011",
--  "11111111111000111001110101100110001011100001110000111101100000000011101001110010",
--  "11111111110001110011110111110010000100111101100010000101111100011111000000010110",
--  "11111111100011101000100001111001101000001110000101110111110101101111000100101100",
--  "11111111000111010100001100111101111111100011000100011011100110000011000001111100",
--  "11111110001110110100111101001101110011100001101011101110001010100100010101010001",
--  "11111100011110011011111100011100000010110110101110001101110111111110101000101010",
--  "11111000111111111110101000100101011011011010100101100111000110011111000001101101",
--  "11110010001100001101010101111100110100010011000100100001001100000011100111101101",
--  "11100101001000000101110011110000101111000101100001000110001000101011001101011110",
--  "11001101000100101110101001011110000011101110001011101101010011001100000000010010",
--  "10100100010001110100110011000000011011111010000110011101101111000001001110111101",
--  "01101001011010110110111000110010001110001100011111010000101011100001000001011111",
--  "00101011011010010100110101111010011111111111111010010010110111010010110011101011",
--  "00000111010111001000101101010111110011001110111101101111110010000010100110000001",
--  "00000000001101100011000100010011010000000010100011011010110111100011110001010010",
--  "00000000000000000000101101111000101111011000011101110001001111101000111110101111",
--  "00000000000000000000000000000000000000001000001110011001001110111101111100000110");





-------------------------------------------------------------------------------
-- ------------------------
-------------------------------------------------------------------------------

--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--use ieee.numeric_std.all;
--use ieee.math_real.all;


----XXX TODO: Maybe split up the ROM into smaller tables. Then access should be
----cheaper and simpler. Use then a distributed RAM. This RAM can also be shared
----with other modules.
----Currently no memory LUTs are used which impacts performance and area usage


--entity ber_eval is
--  generic (
--    MAX_PREC : integer := 79;
--    CONST_K  : integer := 253;
--    MAX_X    : integer := 10
--    );
--  port (
--    clk : in std_logic;

--    --Fifo interface to get randomness
--    rand_rd_en : out std_logic;
--    rand_din   : in  std_logic;
--    rand_empty : in  std_logic;
--    rand_valid : in  std_logic;

--    fifo_ber_empty : in  std_logic;
--    fifo_ber_rd_en : out std_logic;
--    fifo_ber_valid : in  std_logic;
--    fifo_ber_in    : in  std_logic_vector(integer(ceil(log2(real((CONST_K-1)*((CONST_K-1)+2*CONST_K*MAX_X)))))-1 downto 0);
--    fifo_z_empty   : in  std_logic;
--    fifo_z_rd_en   : out std_logic;
--    fifo_z_valid   : in  std_logic;
--    fifo_z_in      : in  std_logic_vector(integer(ceil(log2(real((CONST_K)*(MAX_X)+CONST_K-1))))-1 downto 0);

--    z_dout  : out std_logic_vector(integer(ceil(log2(real((CONST_K)*(MAX_X)+CONST_K-1))))-1 downto 0) := (others => '0');
--    z_full  : in  std_logic;
--    z_wr_en : out std_logic
--    );
--end ber_eval;

--architecture Behavioral of ber_eval is

--  constant MAX_BER : integer := fifo_ber_in'length;
--  constant MAX_Z   : integer := fifo_z_in'length;


--  type bernoulli_vals_type is array (0 to MAX_BER) of std_logic_vector(MAX_PREC-1 downto 0);
--  constant bernoulli_vals : bernoulli_vals_type := (
--    "1111111111111111010010100101001001111000111011101000010110111000100011100111001",
--    "1111111111111110100101001010010101110010110010111110001000001111101010001011001",
--    "1111111111111101001010010100110011101001010100011011000010011000101101001101010",
--    "1111111111111010010100101010000111100001011111111010001100011110110011011100101",
--    "1111111111110100101001010110001111111110000101001100111100010101001000111101000",
--    "1111111111101001010010110100100011100101101000111101100011001100001100001101111",
--    "1111111111010010100110001001010101011010010100100011100101110111011010000011110",
--    "1111111110100101001110010011100000111001111010011010111111000110000100010110001",
--    "1111111101001010100100101010000011010010101001000100100110001100100111111001010",
--    "1111111010010101101001011101010101111100100110001110011011001100000010011100011",
--    "1111110100101101010011001000111000011001001011110101100010011111001110011000001",
--    "1111101001100010100100010101010011011110101000010001110110100011111011110100011",
--    "1111010011100100101010011100110101011010010011100110000110010100001111111100010",
--    "1110101001000100101011111110111001011010100011110000101110010101101001111101100",
--    "1101011001100001101001000000110110101101000101010101101011100111110100100011010",
--    "1011001110000111011000111000010010011000110111100110010010101000110111001100011",
--    "0111110111100110100111001100010110001010010100000000111000111100010100010101001",
--    "0011110111101011000001001101011011111100000010000000111011000000001101110001011",
--    "0000111011111001110110000001000001010110111001011111101000111101010001010011010",
--    "0000000011100000010001110111011111001111101001011100011001101110100011110100100",
--    "0000000000000000110001000111110100100101100111110000111101011011111010100001100",
--    "0000000000000000000000000000000010010110110011111101111011001001010100100110000");

--  --"0000000000000000000000000000000000000000000000000000000000000000010110001101100");

--  signal ber_val : std_logic_vector(MAX_BER-1 downto 0):=(others => '0');
--  signal z_val   : std_logic_vector(MAX_Z-1 downto 0):=(others => '0');


--  signal z_val_out  : std_logic_vector(MAX_Z-1 downto 0):=(others => '0');
--  signal z_val_free : std_logic := '1';

--  signal bernoulli_line : std_logic_vector(MAX_PREC-1 downto 0):=(others => '0');
--  signal counter_exp    : integer range 0 to MAX_BER-1  := 0;
--  signal counter_ber    : integer range 0 to MAX_PREC-1 := 0;

--  type   eg_state is (IDLE, WAIT_RAND, WAIT_RAND2, STORE, BERNOULLI, REJECTION, FIN, WAIT_RAND_AVAIL);
--  signal state_reg : eg_state := IDLE;

--  signal read_once : std_logic := '1';

--  signal bernoulli_bit     : std_logic                    := '1';
--  signal bernoulli_bit_std : std_logic_vector(0 downto 0) := "0";

--  signal next_one          : integer range -1 to MAX_BER-1 := 0;
--  signal rand_rd_en_intern : std_logic                     := '0';

--  signal sample_counter : integer := 0;
--begin




--  process (ber_val, counter_exp)
--  begin  -- process
--    next_one <= -1;
--    for i in 0 to fifo_ber_in'length-1 loop
--      if ber_val(i) = '1' and i <= counter_exp then
--        next_one <= i;
--      end if;
--    end loop;  -- i
--  end process;

--  bernoulli_bit <= bernoulli_line(counter_ber);
--  --bernoulli_bit_std <=std_logic_vector( resize(unsigned(bernoulli_line) srl counter_ber,1));
--  --bernoulli_bit <= bernoulli_bit_std(0);

--  fifo_ber_rd_en <= '1' when (fifo_ber_empty = '0' and fifo_z_empty = '0' and state_reg = IDLE) else '0';
--  fifo_z_rd_en   <= '1' when (fifo_ber_empty = '0' and fifo_z_empty = '0' and state_reg = IDLE) else '0';

--  rand_rd_en <= '1' when (state_reg = BERNOULLI and next_one /= -1 and rand_empty = '0') else rand_rd_en_intern;


--  process(clk)
--  begin  -- process c
--    if rising_edge(clk) then

--      if next_one >= 0 then
--        bernoulli_line <= bernoulli_vals(next_one);
--      end if;


--      z_wr_en           <= '0';
--      --fifo_ber_rd_en <= '0';
--      --fifo_z_rd_en   <= '0';
--      rand_rd_en_intern <= '0';

--      --Final buffer
--      if z_full = '0' and z_val_free = '0' then
--        z_dout         <= z_val_out;
--        z_wr_en        <= '1';
--        z_val_free     <= '1';
--        sample_counter <= sample_counter+1;
--      end if;


--      case state_reg is
--        when IDLE =>
--          if fifo_ber_empty = '0' and fifo_z_empty = '0' then
--            --fifo_ber_rd_en <= '1';
--            --fifo_z_rd_en   <= '1';
--            --state_reg      <= WAIT_CYCLE;
--            state_reg <= STORE;
--          end if;

--          -- when WAIT_CYCLE =>
--          --   state_reg <= STORE;


--        when STORE =>
--          --Store both values in a register
--          if fifo_z_valid = '1' and fifo_ber_valid = '1' then
--            ber_val     <= fifo_ber_in;
--            z_val       <= fifo_z_in;
--            counter_exp <= MAX_BER-1;
--            state_reg   <= BERNOULLI;
--            z_wr_en     <= '0';
--          else
--            state_reg <= IDLE;
--          end if;


--        when BERNOULLI =>
--          if rand_empty = '0' then
--            if next_one = -1 then
--              --If there is no more onw, then we are finished
--              state_reg <= FIN;
--            else
--              --A one has been found
--              counter_exp <= next_one;
--              --state_reg         <= WAIT_RAND;
--              state_reg   <= REJECTION;
--              --rand_rd_en_intern <= '1';
--              counter_ber <= MAX_PREC-1;
--            end if;
--          end if;


--          --when BERNOULLI =>
--          --  --Do the rejection sampling
--          --  --There should be randomness available
--          --  if rand_empty = '0' then
--          --    --Whole poly has been checked -> Finished
--          --    --See if a one bit is set, then do rejection sampling
--          --    if ber_val(counter_exp) = '1' then
--          --      rand_rd_en  <= '1';
--          --      state_reg   <= WAIT_RAND;
--          --      counter_ber <= MAX_PREC-1;
--          --    else
--          --      --Some more logic, to search for zer
--          --      if counter_exp > 2 then
--          --        if ber_val(counter_exp-1) = '0' then
--          --          counter_exp <= counter_exp-2;
--          --        else
--          --          counter_exp <= counter_exp-1;
--          --          rand_rd_en  <= '1';
--          --          state_reg   <= WAIT_RAND;
--          --          counter_ber <= MAX_PREC-1;
--          --        end if;
--          --      else
--          --        if counter_exp > 0 then
--          --          counter_exp <= counter_exp-1;
--          --        elsif counter_exp = 0 then
--          --          --The last bit is not one, we can accept
--          --          state_reg <= FIN;
--          --        end if;
--          --      end if;
--          --    end if;
--          --  end if;


--        when WAIT_RAND =>
--          state_reg <= REJECTION;

--        when REJECTION =>
--          if rand_valid = '1' then
--            if (bernoulli_bit = '1' and rand_din = '1') or (bernoulli_line(counter_ber) = '0' and rand_din = '0') then
--              --Nothing happened - no decision made
--              counter_ber <= counter_ber-1;

--              if rand_empty = '1' then
--                state_reg <= WAIT_RAND_AVAIL;
--              else
--                state_reg         <= WAIT_RAND2;
--                rand_rd_en_intern <= '1';
--              end if;

--            elsif bernoulli_bit = '1' and rand_din = '0' then
--              --smaller = accept this line. See next lines
--              state_reg <= BERNOULLI;
--              if counter_exp = 0 then
--                state_reg <= FIN;
--              else
--                counter_exp <= counter_exp-1;
--              end if;
--            elsif bernoulli_bit = '0' and rand_din = '1' then
--              --greater = reject
--              state_reg <= IDLE;
--            end if;
--          end if;

--        when WAIT_RAND_AVAIL =>
--          if rand_empty = '0' then
--            state_reg         <= WAIT_RAND2;
--            rand_rd_en_intern <= '1';
--          end if;

--        when WAIT_RAND2 =>
--          state_reg <= REJECTION;

--        when FIN =>
--          if z_val_free = '1' then
--            state_reg  <= IDLE;
--            z_val_out  <= z_val;
--            z_val_free <= '0';
--          end if;


--      end case;
--    end if;
--  end process;


--end Behavioral;

