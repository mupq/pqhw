--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/

--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:58:31 03/01/2014
-- Design Name:   
-- Module Name:   C:/Users/thomas/SHA/Projekte/BLISS/code/bliss_arithmetic/lattice_processor/verification_finalization_tb.vhd
-- Project Name:  lattice_processor
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: verification_finalization
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

entity verification_finalization_tb is
  generic (
    MODULUS_P_BLISS : unsigned := to_unsigned(24, 5);
    PRIME_P         : unsigned := to_unsigned(12289, 14);
    ZETA            : unsigned := to_unsigned(6145, 13);
    D_BLISS         : integer  := 10
    );
  port (
    error_happened_out    : out std_logic := '0';
    end_of_simulation_out : out std_logic := '0'
    );

end verification_finalization_tb;

architecture behavior of verification_finalization_tb is
  signal end_of_simulation : std_logic := '0';
  signal error_happened    : std_logic := '0';


  signal clk      : std_logic;
  signal az1_data : std_logic_vector(PRIME_P'length-1 downto 0)         := (others => '0');
  signal c_data   : std_logic_vector(0 downto 0)                        := "0";
  signal z2_data  : std_logic_vector(4 downto 0)                        := (others => '0');
  signal coeff_we : std_logic                                           := '0';
  signal u_out    : std_logic_vector(MODULUS_P_BLISS'length-1 downto 0) := (others => '0');
  signal u_wr_en  : std_logic                                           := '0';


  -- Clock period definitions
  constant clk_period : time := 10 ns;

  type ram_type is array (0 to 512-1) of integer;

  signal az1 : ram_type := (801, 2228, 4750, 5266, 10684, 683, 8114, 1667, 8115, 2955, 4440, 7178, 10196, 6621, 8571, 2797, 1588, 6394, 1076, 3127, 9288, 3322, 3523, 9767, 191, 6861, 11701, 2365, 5749, 10998, 6120, 1200, 1765, 2792, 3593, 6567, 9859, 6785, 790, 11917, 5703, 890, 1918, 8832, 6313, 10372, 11837, 7564, 6402, 158, 1833, 11773, 2636, 4674, 748, 12207, 11245, 11354, 10461, 1204, 8504, 7933, 945, 4012, 7193, 9320, 10411, 3696, 2239, 11751, 9205, 7084, 7761, 4144, 5502, 4877, 12224, 9224, 11275, 11707, 12033, 4170, 1652, 4584, 4516, 3625, 6698, 1226, 7321, 1120, 7800, 7780, 3133, 5678, 11342, 810, 12255, 9491, 5875, 9105, 10370, 9317, 11678, 2479, 10633, 2224, 6606, 9114, 8440, 1936, 9708, 6840, 12196, 10364, 7427, 8583, 10028, 10787, 8002, 7040, 646, 5509, 7397, 11413, 9335, 9402, 4911, 10486, 10075, 8959, 2991, 1412, 10625, 1576, 153, 2367, 3574, 2762, 5277, 6750, 1549, 10400, 2076, 569, 12036, 8169, 4725, 6755, 6547, 2882, 1458, 10262, 8211, 5286, 9525, 6439, 9318, 10182, 5791, 7732, 9318, 6189, 1288, 3599, 1423, 2646, 8330, 5900, 7185, 5636, 6922, 10140, 10027, 11825, 10500, 2104, 596, 10419, 1999, 10212, 10728, 11480, 7719, 2940, 1787, 5435, 9027, 1509, 2081, 3687, 1317, 4288, 11643, 666, 1246, 10254, 6901, 8616, 4144, 11002, 2145, 438, 1186, 6044, 938, 3223, 6958, 4369, 1591, 3680, 2444, 3526, 2141, 10366, 218, 4819, 3653, 1550, 6620, 5127, 10306, 8195, 11046, 10818, 5413, 12224, 3489, 203, 10000, 1278, 8250, 5453, 2758, 9856, 9097, 6089, 8888, 98, 8483, 11603, 7727, 1355, 5917, 741, 6895, 10320, 4176, 737, 2160, 8562, 7358, 6899, 9849, 8846, 1805, 7282, 6927, 7218, 906, 9730, 7526, 11378, 3262, 9188, 3325, 3792, 9728, 7507, 11172, 8167, 2507, 7751, 2725, 2492, 3752, 2877, 5849, 11995, 10635, 8671, 10316, 12149, 9348, 3593, 11151, 8996, 11908, 11607, 10356, 10103, 5475, 3628, 11750, 8125, 7334, 12052, 3098, 8637, 180, 7464, 3226, 9676, 3937, 188, 2478, 9562, 2803, 2378, 95, 10681, 271, 6325, 6801, 11440, 5938, 6143, 11719, 7743, 5669, 9191, 958, 4144, 6520, 5873, 10540, 1860, 1606, 11369, 1091, 379, 12263, 5829, 7713, 6421, 4466, 4503, 3316, 11238, 3721, 9306, 8033, 3957, 7793, 5810, 1084, 8820, 9912, 9729, 2872, 5117, 4866, 3227, 3571, 9116, 5494, 11180, 5353, 11889, 970, 7843, 1240, 11210, 6323, 7644, 6968, 11089, 5570, 3265, 9388, 6610, 9317, 9018, 7993, 5496, 5128, 4762, 3811, 11228, 2654, 7983, 5640, 8190, 8532, 7333, 4699, 6135, 9776, 4804, 10464, 8542, 3332, 12247, 5041, 1365, 11044, 9986, 6016, 7271, 2191, 2555, 11537, 2108, 6610, 3292, 3828, 1034, 6505, 4528, 2935, 11019, 10226, 265, 1773, 11393, 10173, 4386, 12099, 3271, 1708, 6994, 11078, 9171, 1162, 1094, 8024, 8505, 6885, 9188, 7376, 2557, 2849, 1264, 1287, 5765, 2090, 2542, 744, 6848, 6250, 386, 12006, 3362, 38, 489, 1200, 9116, 4299, 3570, 1633, 5126, 7207, 12077, 8027, 2926, 9747, 5195, 775, 1805, 4486, 7338, 6292, 10767, 7684, 4689, 6555, 8645, 11861, 2593, 5591, 10557, 1591, 9144, 5374, 6848, 1800, 12087, 1043, 8799, 3895, 5179, 4560, 12101, 7508, 10184, 1707, 621, 4395, 439, 10641, 8795, 9529, 7636, 2732, 1656, 3972, 5655, 2853, 6803, 2809, 8122, 10716, 6084, 272, 6946, 11457, 1366, 3629, 11514, 6259, 2151, 2367, 1208);

  signal c : ram_type := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);

 signal z2 : ram_type := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0);

  signal result : ram_type := (-11, 2, 5, 5, 10, -11, 8, -10, -4, -9, 4, 7, 10, -6, -4, -10, 1, 6, 1, -8, 9, 3, -9, -3, 12, -5, -1, -10, -6, 11, 6, 1, -11, 3, -9, -6, -2, -5, 1, 0, -7, 1, 2, 9, -6, 10, 0, 7, 6, 0, -10, 0, 3, 5, 1, 0, -1, 11, -2, 1, 8, 8, -11, 4, -5, 9, -2, 4, -9, -1, 9, 6, -5, 4, 5, -7, 12, 9, -1, -1, 0, 4, 2, 5, 4, -9, 7, 1, -5, 1, 8, 8, -9, -7, 11, 1, 0, -3, -6, -3, 11, -3, 11, -10, -2, 2, 6, 9, 8, 2, 10, 7, 12, 10, -5, -4, 9, -1, 8, 7, 0, -7, -5, -1, 9, 9, -7, 10, -2, 9, -9, 1, -2, 1, 12, -10, 4, 3, -7, -6, -10, 11, 2, 12, 12, -4, -7, -6, -6, 3, 1, 10, -4, 5, -3, -5, 9, 10, -6, 7, 9, -6, 1, -8, -11, -9, 8, 6, -5, 5, 7, 10, -2, -1, 10, 2, 1, -2, -10, 10, 11, 11, -5, 3, -10, -6, -3, -10, 2, -8, -11, 4, -1, 1, 1, 10, -5, 8, 4, -1, -10, 1, 1, 5, 1, -9, 7, -8, -10, 4, 3, 3, -10, 10, 0, -8, -8, 2, 7, -7, 10, -4, 11, 10, -6, 12, -9, 0, 9, 1, 8, -7, 3, 10, -3, -6, 9, 0, -4, -1, -4, -11, -6, -11, -5, 10, 4, 12, 2, 8, 7, -5, 10, 9, -10, 7, -5, 7, -11, 10, 7, 11, 3, 9, -8, 4, 10, 8, 11, -4, -9, -5, -10, 2, 4, -9, -7, 0, -2, -4, 10, 0, -3, -8, 11, 9, 12, -1, 10, -2, -7, 3, 11, -4, 7, 12, 3, -4, 0, 7, 3, 10, -8, 0, 2, 9, -9, 3, -11, -1, 12, -6, -5, 11, 6, -6, 0, -5, -7, -3, 1, 4, 6, -6, 10, 2, 1, 12, -11, 12, 0, -6, -4, -6, 5, -8, -9, 11, -8, 9, -4, -8, -4, 6, 1, -3, 10, -3, 3, -7, 5, -9, -9, 9, 5, 11, -7, -1, 1, -4, 1, 11, -6, 8, 7, -1, 6, -9, 9, 7, -3, -3, -4, 6, 5, 5, -8, 11, 3, -4, 5, 8, 8, -4, -7, -6, 9, 5, 10, 8, 3, 0, -7, -11, 11, 10, 6, -5, -10, -9, -1, 2, 6, 3, 4, 1, -6, 5, -9, -1, 10, 12, -10, -1, -2, 4, 0, -9, 2, 7, 11, -3, 1, 1, 8, -4, 7, 9, 7, -10, -9, 1, -10, -6, 2, 3, 1, 6, 6, 0, 12, 3, 0, -11, 1, 9, -8, 4, -10, 5, -5, 0, -4, 3, -2, -7, -11, -11, 4, 7, -6, -1, 8, -7, -6, -3, 0, -10, -7, 10, -11, 9, 5, 7, 2, 0, 1, -4, -8, -7, 5, 0, 7, 10, -10, -11, -8, -11, -1, -3, -3, 7, 3, 2, 4, -6, -10, -5, -9, 8, 10, 6, 0, 7, -1, 1, -8, 11, -6, -10, -9, 1);

  signal counter : integer := 0;

--signal az1 : ram_type := (3143,8726,6251,11273,7202,11610,2469,1640,2799,6726,2096,11224,8492,12075,2030,7659,1766,4050,3170,4974,198,5861,8641,5952,1054,9872,1865,8784,4319,1993,668,4970,4505,8245,8817,3358,11558,8826,11410,9259,5467,5125,2383,7807,6820,10726,1903,9686,1053,11436,11223,2958,5272,7348,9506,3745,10104,8944,6495,1953,8213,6154,1448,1,5422,1621,9088,9260,4952,9115,7254,5134,3772,1599,2613,11759,1972,11155,3300,10470,420,5951,9001,11746,10628,3885,1625,12174,11471,7730,10817,12150,5785,39,1577,7039,2110,1880,4300,7543,2043,1026,10856,2096,7281,715,11550,4603,11153,7917,2890,1728,11648,12280,5847,8035,5619,7145,10081,9646,3877,1166,3,8280,1315,2507,10913,3532,10856,11281,9455,4048,11871,4105,10341,909,9858,2485,2955,12006,11235,4031,10062,4043,7150,8798,7047,8698,1848,10143,11461,405,7657,3964,1553,5893,7716,4559,3913,2082,3454,334,613,7018,6859,897,3463,729,2944,5373,3963,4564,10849,2583,11037,6968,10548,3479,108,4691,2418,5507,9852,11410,756,7135,5593,4210,3346,10905,6711,6492,3400,6107,515,2360,2139,804,12204,9214,2418,12210,9195,6851,7884,11509,4032,249,652,11003,7751,6069,5201,431,6304,3418,11962,188,11812,3530,5849,4670,4414,10325,10920,231,4430,2877,1945,3052,3736,10649,978,11950,3266,295,10772,8916,2375,6417,4251,279,4664,3219,8380,3483,425,3862,1731,1420,6885,2601,7046,3261,3817,7810,4386,615,139,7084,10818,2836,858,8581,8876,10180,8912,11815,4347,4181,11971,8420,752,11286,4793,10778,3715,9858,11421,10588,2999,7183,7583,1299,5502,3437,2854,4335,6400,4307,227,6418,7030,10769,2743,2094,550,9234,1743,112,2805,11461,6174,8787,7989,9165,3320,8335,5071,8864,10432,4155,7877,9728,11977,1015,1496,4079,6373,10252,10214,12235,3109,9831,8562,8981,281,2490,11119,6869,3328,2378,5817,11402,5356,6545,7706,9421,12143,5601,11451,4486,3953,12257,5154,11126,799,8294,4598,75,405,2885,2581,4044,11710,10705,8776,8812,4396,5023,3141,10418,4784,9798,5675,4667,8302,10595,5705,721,4826,3138,5165,7317,4320,4156,1773,11950,5138,1653,8897,10444,6717,11462,12016,8468,4743,5167,3026,4662,2507,3925,1909,1356,4821,1261,7739,9264,11465,6379,4702,7409,1255,4205,11644,8084,10711,6035,5164,7155,4175,7318,5077,9817,990,5961,4177,377,3064,115,8538,9205,6524,5189,2913,9721,10533,6709,5058,12269,8896,2624,1765,10131,7415,9319,5478,4822,5879,58,7183,9147,5727,6877,5339,9127,10514,11108,11533,9573,481,9654,2299,5569,4543,1737,4117,4984,4427,2736,9839,8950,83,4217,7627,8468,8544,1148,5471,2830,10734,8279,10759,8690,8883,1876,7440,5958,1237,10770,8633,9539,1251,4776,6048,6759,10572,10424,7117,9289,6827,10681,8414,5205,2963,11785,10052,3585,10869,7325,2328,3593,5211,11779,7647,3793,9514,1567,5688,350,10683,3647);


  --signal c : ram_type := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0);

  --signal z1 : ram_type := (263,232,-361,154,-29,-55,15,380,-474,-243,-22,-494,-258,-110,640,47,-90,211,-31,136,-133,-9,102,179,199,302,428,-146,176,-206,-172,-14,-497,-341,172,126,151,51,46,198,138,205,181,-5,-120,297,442,131,131,148,-234,-140,-45,-285,170,135,181,-425,-47,130,-399,31,-39,-167,455,-243,-312,-105,220,229,337,-18,-176,-69,104,-139,145,-13,-147,-10,145,-5,-468,274,59,-259,-144,118,123,267,25,324,187,-212,320,-217,-108,163,71,-90,59,-191,117,309,329,-86,234,166,66,140,-247,-140,-187,-222,-154,-260,16,-130,-43,358,-80,-287,228,-2,102,-135,-144,362,-91,-198,-79,75,141,-80,256,290,18,96,-351,118,545,121,-216,-402,133,83,-111,-106,-24,-181,419,-259,188,94,-10,41,373,10,170,-250,-629,58,140,403,-142,-125,62,-367,370,-207,181,-179,67,37,-70,16,208,-255,141,-188,298,169,-24,107,-91,-97,-6,295,-128,-78,-207,110,-171,347,7,-16,37,-77,-162,-70,-233,-134,-5,-226,128,351,-155,-167,-32,104,24,72,74,-49,-98,-47,208,150,-314,-103,-120,122,420,48,-268,-43,-99,154,197,121,-554,-199,179,-125,-171,79,-503,-193,-381,160,59,-104,230,99,151,-382,-231,202,-39,-12,-25,375,243,393,-215,19,-114,164,217,-300,112,70,217,-89,291,-159,89,-14,207,-392,454,-75,-133,118,-280,138,464,-377,476,-72,413,85,-351,-211,-95,95,378,23,336,273,-233,18,-349,259,73,383,443,98,193,-298,186,-43,-38,-47,299,-71,-38,-170,-120,-380,-219,-27,183,-151,171,224,548,164,-173,-302,-502,-598,-142,-515,-34,-151,-25,-188,-53,-154,7,5,87,-211,-262,-64,-536,249,-458,164,189,-24,-199,-58,99,238,33,315,115,131,119,-112,-121,508,366,-301,-190,-441,176,304,-115,147,49,16,-310,117,14,74,-127,-296,367,58,288,-1,-96,-207,-54,-47,-39,-197,633,-121,149,-6,148,332,-398,-165,-293,391,-141,-16,-75,-282,0,147,-220,-313,120,-55,46,16,59,145,-412,-278,184,141,-84,239,240,-300,-107,319,-199,-83,62,373,365,-480,-224,32,311,-162,-381,470,-14,69,76,3,223,9,-13,-271,123,-88,-113,-150,-8,-280,196,-91,10,-273,165,52,175,-321,-157,-65,260,-159,-197,205,73,-18,-298,143,265,-186,-263,170,535,-16,-475,182,186,-14,400,-89,-23,-122,139,-274,-394,-93,-186,-134,97,195,160,-184,112,147,-296,-204,57,105,-474,85,445,-51,143,-58,-40,91,84,111,95,-11,366,111,-190,100,399,215,-31,-21,-110,-302,-49,150);

    
  --signal z2 : ram_type := (0,-1,0,0,0,1,1,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,-1,-1,-1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,-1,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,-1,1,0,-1,0,-1,0,0,-1,0,0,0,0,0,0,0,1,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,-1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,0,0,0,1,-1,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,0,0,0,-1,1,1,-1);

 --signalresult : ram_type :=(-9,8,-6,-1,7,12,-9,2,-9,6,2,11,8,0,2,7,-10,4,3,5,0,-6,-3,6,1,10,-10,9,-8,-10,1,5,-7,8,-4,3,11,8,11,9,-7,-7,-10,-4,7,11,-10,-3,-11,11,-1,3,5,7,9,-9,9,9,-6,-10,-4,6,1,12,5,-10,9,9,5,-3,7,5,4,-10,-9,-1,2,-1,3,11,0,-6,-3,11,10,-8,-10,12,-1,8,-1,12,-6,12,-10,-5,2,2,4,-5,-10,1,11,2,-5,-11,11,-7,-1,-4,3,1,11,12,-6,-4,-7,-5,-2,9,-8,1,12,8,-11,-10,-1,-9,11,-1,-3,4,-1,-8,-2,-11,10,-9,-9,0,-1,-8,10,-8,7,9,-5,8,2,-2,-1,-11,-5,4,1,5,7,-7,-8,2,3,0,-11,7,-5,-11,-9,-11,3,-7,-8,5,-1,-10,-1,7,10,-9,0,-7,2,-7,10,11,1,-5,-6,4,3,-1,-5,6,3,6,-11,3,-10,-11,12,9,2,12,-3,7,8,-1,4,-11,1,-1,-5,-6,-7,12,6,3,12,0,-1,3,-6,5,4,-2,11,12,4,-9,-10,3,3,-2,1,12,3,12,10,9,-10,-6,-8,-11,-7,-9,8,-8,12,4,-10,1,-5,-9,7,-9,-8,8,4,-11,12,7,10,3,1,-4,9,10,9,-1,-7,-8,-1,8,0,11,-7,10,-8,10,-1,-2,-9,-5,7,-10,6,-9,2,-8,6,-8,12,6,7,-1,-9,2,1,9,-11,0,-9,-1,6,-3,-4,-3,3,-4,-7,-3,10,-8,-5,10,0,-11,2,4,-6,10,10,0,-9,-2,8,-3,12,2,-1,-5,3,2,-6,11,5,-5,7,-3,11,-7,-1,4,-8,0,5,11,-11,8,4,12,12,-9,-9,4,11,-1,9,9,4,-7,-9,10,5,10,-6,-7,8,10,-6,-11,4,3,-7,-5,4,4,-11,0,5,-10,-3,10,-5,11,11,8,-8,-7,3,5,-10,-8,-10,1,-7,-10,-5,9,-1,-6,5,-5,-10,-8,11,8,-1,-6,5,-5,-8,7,-7,-3,1,6,-8,12,3,12,8,-3,6,-7,-9,-2,-2,-6,5,0,8,3,-10,-2,-5,-3,5,5,-6,0,-5,-3,-7,-5,-7,-3,10,11,-1,-2,-11,10,-10,-7,-8,-10,-8,5,-8,3,-2,9,12,-8,-5,8,8,1,-7,3,10,-4,-2,8,-3,2,7,6,-11,11,-4,-3,-11,5,6,-6,10,10,-5,-3,-5,-2,8,-7,-9,0,10,-9,-1,-5,-10,-8,-7,-1,-5,-8,9,-10,5,1,-1,-9);


    
begin
  verification_finalization_1 : entity work.verification_finalization
    generic map (
      MODULUS_P_BLISS => MODULUS_P_BLISS,
      PRIME_P         => PRIME_P,
      ZETA            => ZETA,
      D_BLISS         => D_BLISS)
    port map (
      clk      => clk,
      az1_data => az1_data,
      c_data   => c_data,
      z2_data  => z2_data,
      coeff_we => coeff_we,
      u_out    => u_out,
      u_wr_en  => u_wr_en);


  -- Clock process definitions
  clk_process : process
  begin
    clk <= '0';
    wait for clk_period/2;
    clk <= '1';
    wait for clk_period/2;
  end process;


  process(clk)
  begin  -- process
    if rising_edge(clk) then
      if u_wr_en = '1' then
        if u_out /= std_logic_vector(to_signed(result(counter), u_out'length)) then
          error_happened <= '1';
        end if;
        counter <= counter+1;
      end if;
    end if;
  end process;

  -- Stimulus process
  stim_proc : process
  begin
    -- hold reset state for 100 ns.
    wait for 100 ns;

    for i in 0 to 511 loop
      az1_data <= std_logic_vector(to_unsigned(az1(i), az1_data'length));
      c_data   <= std_logic_vector(to_unsigned(c(i), c_data'length));
      z2_data  <= std_logic_vector(to_signed(z2(i), z2_data'length));
      coeff_we <= '1';
      wait for clk_period;
    end loop;  -- i
    coeff_we <= '0';


    wait for clk_period*1000;



    if error_happened = '1' then
      report "ERROR";
    else
      report "OK";
    end if;

    end_of_simulation <= '1';
    wait;
    
  end process;

end;
