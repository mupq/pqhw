`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VsinksLpJWI1tuaOI7h8aSORfn/+DW4FgGWyEDOqHNlVivfJQf+MdvTR8ppGqPOJph04UfQew3Tt
9UcXkhvcCQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+q7wFKp4PHZ99AOUXOfirVj8vjzVgTcROZi67zAuw/5nj1fUNd8IrtLm017VkcF7WHeCEaKQOit
7blqlCcFByKHzQZW2lCOHhJ9lEeJxJj967u6BCbISZhlKVikQBA8fKRVVZn0WvcMZn77lmVL7JTc
D8KSr6wy9yJwkkV+ppg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W2UVrope1p5WH2sS/2M7d2v+U87r5bZ1kcQCK80etZcsJN7glyuCz7NAnFVTiQhwq2JxwCBoVOEf
8BNELEM0HOxMWOFqPzWztADNCxArYYKM7CGbUSiNCCD4bdpKHBPHGPYVs4ePAKJGoVYgB8JAz9cG
Aa8RBN5Qx71Y9FxO58FCXPFCc6UTW26PNiGdlVOGG182Blnfw2zmLnNc/DXqiUa/NQKsDHrDwxHR
XPsvWVIUh6+IU5hYZZJwEqWBcm4bj4I16etHiYIe+EPeftbKa6UcdBWIzYmW0Bz2WOn7tCADIUpM
PifKVu5RzyoJjNiGbp9Z3S9dpTJynoDuBvID9w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h6rZV2rYxkx1Ra2F0CM6473N9Mzbp8xIWRu0//VbQefhQbOMXtTVTxhCItdVdR4EfFsRZVI7+nt7
9KJ7Um1ycu0Gx2wyjgWOmLlY2v62OYdx4w7yId4HA35a4yo2J6/kKJYlM00NmVziarFDB7al9/de
EwEjHKg7DQl0oyrlbvw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bv4R6oBTTV/Ekm8xZ5sZQat0BLfpO8TeLbF1+Xcd6TrfhzW5K3nQ80+HK8qvK6o6zcyKypall82o
bEISra9NsvpO17A/MNcMY8Jvt4J+nlPv2hZqLiR4f/Tau55kV3j+FopH6wzcicrl672uRYGgNBB6
wPEhmpqGHrIloK11m124q5xZEHCZmz+16YsroAgM8nfdm7r8dBytwyF5338RSeK8MlbvBR8kYUFx
f30JLB2q9/nlc57jD1fhdTsLKIaxFI6L/hh4l+vWb3d2FG0fW1mQJnB0omomUYLkfezFp/WkmP+X
JoEz3xpGC/PExNVEwJnGKnFX4uSp2hZRTx46Wg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LSNZAyyvsFlTnG6tGAEv7pRHmgtMyJkEsbP6DfPx7YLChIw7VTeSUXKqKiSxcdFMzbEH6PVN5OXU
TOzOe4LQSB4VrDpMHU1iWuuQK5hU6V+wT9+NKx1cCF2+4zfr2alMgIb9PGOgArGsXYvJBEEKTH7v
SQ2wXjEs8OBK/1ScP8hDVuAAHMTRDlfU4a9W50nqxIHdJOzL5EPbQa2W1W3sEyJ51s0yVcASBMwH
b+rBsOhU6NgQuKQ6DQj9VNNr7myYq7PN/TIdYKSzLOuFMm7bG7gu7rUs7LtIxQeSI2Z4K70PKGJF
OVJKu6LUG9jJJXt7UlnU74Siw0CA/SX0KpbOOw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17440)
`protect data_block
IP/Wr3Q3IiSmAivHcrmPxdvvGQKkce6vuS8vhwWgV1bTcffY/oeMmcaaWVxhJAy6QJcSq6oBstOm
WAwr2KZi0tw3PBF1gIASoQPg1TAJoJB6PITDwNuALCsmYfVNdxxk5EoTYYhvJrx2p6E+Tq/dlvas
K5y5jtTZX53zkcT1en/RlLLPkyoplKTRMFxkoPzzUjr2AjVoygDEyx0w3ZXPuhTzATqg6GsGguZu
vlA/oir9tmW25m5axXr+6YGVdrmLaHs+JUPq3u/AgsbYD2rfwbkeVasxKioa56suQROAHZvKt8T9
6RyGpy71SzN1jMYm1ywciVr925xdsqsZIKwT2LSB0nbgd7hHD0hlOHDG5O1HrtEYqpYzRPO3GISM
Ff1ED3CThyWY/i2Nk8VL23ar5vyCePdCHB53IfC/QX8kWClqeJ/FmrSy7sP1So/pB8AabvWr3Hja
Dudz8XJpBdwN7xV8TWYz/NGo+WIk0/RR5qUc9WJ+Y16ULe8X5FzQqalWuA4IH13j7CoKSxhGACbL
lzp7rLM3P1IByWHw0B3La0NMQ5k1Kz6W9qlzJ2V00q/DSb9Gv6SsgbASgFuY+HgqtxCLOgsLlTvw
c1v2/SufiYv7OFiwvn7FKybWJCukMUTx6na6q62V912i0HCI0azQ1pgPXK2kg6LEYKolpam89LiA
2ITUT7Aq7mEda7trOTo4IxB2wpuWLWMtH6+62S6Qm0mNbNUqQO4SWo2vA1ZvDhNXXLtDtgCTkIAY
Pxe4p1zR+VTGybsyF3+Rx6K2tsz+znlt6btY5qhy5K0olqMUZUthipjS2cs4S//PeGDTcv5581/U
qfXL9Ti9h12GYhf+NY9DBD8sX4aDW1hjgWFVlM/Vlv0Jr+GXCyv9tv64byekFaPrF6ahFdSGy+bv
f5zLGma57rJWo8gTmt+GShwdI9aUhkHStiJ968yhbrGZkfI5YcxbTkNYYAwFhqaq0PFWpxXPxPW9
VGrgab52TqGZ6kawkwJrzKx0lxx1UrwwWNb17xSFDLv5h6XOal2ldjo8950SGBs+mKn5LNK0d1T8
a53X6/+rWNfDc9120PxqcQ75RZ1Ex+BUOAhPlYfQpIspUHtxjm6nGKNYoIaduYwcqXTjIh88IHni
Vw7gbHXFMzGWJETRx7YY9hPGFQLxD1uJEkWfn6kEF9l4Q7f6pn+83Btn0c1MfKjmA6Dn9itgTguL
7brxxlrg9upfvi3IbAiU40aOAOozNgUxhoAl3VajhSghwfCEx8G0whNKxdXAJHZFRUrgg1YXZJRk
5A6BM9PehHZzIsmimmQX58LFl8k/U3snadxfsB2OmW2mJY+BqYML89y3bxy79DLVsfEuchsA9X2v
v3S0lW7xSSEo9Grlw96/XngUdhr13DFEkk+P+HsPgkUKWkF8/REBH8Eg2Qd9f4O3HHIiPHLKd8y7
BbxBj4Xb6/r3t+25fn/KXZ6NvE41ZFCjD1WgQvsZN60nRuxCiIgST29WaHNjOeZd0s76zZsx96uO
4B7RWGjobG6J/MUbkv9Io4NUnOHRhnAMVp24V7A0dqyAh35gjZ4rdmHjCK977IG1+1Uo5Ddtfcd6
MqjPvFSB1d/XdbWpVchGKqle2I8dQsY2rmZiA4dXOARP5e7xpZ8Xt1WfVZq8AZS/6TE0GhIFHqgF
kQA96+V8mHW4tCFwdCPh47Dze7+BmbCnecU0LlmsH/WJxKu+0XO8feUkpSEj3uGikBlm0XitLSfs
y5/rgiR8MewQmhrMMK3F/kS9sRx8CAuY7VFOfPL5sVRJ5T9fNWnU+D/Uqffy38OaR2WH391wfziF
tFubFYGkocGTkGd6zHksfGnPPSZLKRqfpRmbCgjO5qkXuCZKioIXNk8lI76dNwoeO+7blW0pGGcx
NT2BJLn0P2qfx6BZCEFTRILBCn4lwhXUI2XeRkKl8Wa6q8MdcbUx0LhtN5ZmuIbQEclLRPhlRqFR
rD1lVwmMgR9h5AoTb7PWtFjOvQ/Zw6SWwJLr7srPc/GVnUNUM064IpRjHvVZpwUG7bVPZUBdl8h2
u7Px5aDZgHwPumAcziqImpA3qQ30I03WIq13cto0pAj5zGCE310D5wLELrqfUFUcHVWQ/O0pqUH3
ognbE7XKJXVxsb+eZOkVGjVvWh8XCG+jQEWV+ENbZ5rF+XFbyqSYjMWuAJMUFDRX/X0W0XL/IOlN
dHfLYzYuEv5CFz2tHvdNsrkLph0AJ/jVVj9Axro357VjPbYvg68WHnK2Fsc6hjvZqqwG/0Yvn44Y
8QncTKRgZJp+F/gOqhTFUShXVyslcZGP4QZBAzhPuX8RnXx1cjYpIKCE79veMngYGUNuTKyP+8sx
H2H+1xCtwNPQs3UwbSVJA9j/Q6NittfmlbpsrbkhPabmot5g+6Eqh7/PhyudVRHSBsN9IHO9B430
HNGDPzJsfE2ZPkJJz9MuDryw7cYqhZEpwepJxxyihVUsupZaMD0yfeKDIxjCglRRXQidbAQFjQ//
268psMzzasB4stLqyNAFmKuf/SogTDehIbEjAPKE0XrG2RN7SiVr6E1eZpoMr8P4BS764iEnWzIC
vTCJqbHnN040RnlyI+cHrX1PHh+vmSev23HifuSXt1EZWFI/mHfQp1wVZwiYR09ti6uJIrQoFPr+
7oCt/A/ntzYrMiPVn7/HIOMXuewXjWZQsMFH8fsi2piJ+ubln67KW4neCwUMsta8FPg6cEQlXrVD
+l2uxxbi4kTOkvLTn6MEwX/UmmMqKPdnkUsFL3AKpjH/7VP2o9OLOWhQh4wzNS6bejb+MpN7XZGy
IyQZmUccwovhIYk0TcwRtputIU/87TGWLULxDwPW8RlXnFL807tB4jv6vYM9xVutVfgVTRcIoH7L
uANhovEdFMcLDNxio0P+uDuy2jh4r5TKCUh5tWFluHwxKFsjrLvRKZyuCET6wzOXybKzWJBSEZHh
1owEoPKLHKwfSt27JbnOs+n3A3pTqD000Fu/MopoicyMAF2XOSsB8X4gj2wwEHM9eNTLLaHAGJTo
jyjKj2npf05oUuZ2cWkw5v6gVXhg6oGM0Uasw8q5ewN9qLZWPL2q5KtgmomHg5hMtCVQQOgBhntP
3cbW0WG4fALe2Co8NWib+g2QRtL+RlqQxevo+BItSUti/aUrCFHvwt25nTB17nHsBteNElvMyfz/
Z3/PTmW8OeEgW9B7YGfhbzkwJn/IVyIO8zMlNXz2CVOIlhI7H+WNJL8KYZJ1hKyLXxkd5KAOI+KJ
OLVP0pQKxOsgjM4Jm/x5NFgK1lYr+WjO0W24gHBcI0+GzT7QFhnkdsDp1p2/DE1PCrjh/WAul6Ni
7xkzKnVUNmpYdwrTC0VSKXll9yf8Z9FRoTFkcrLnyenqqSD9uDKOkBN1B+uy6864V65NrEoUAJYW
IcM9w3kyXg4tRVSvG565KyG7TsBHSyUFFexK/d90N6HyZP08SuB5wv4fL/RRvXFvCRBXtv/X88h5
IB93nQ6TvVfydEnigCLLvDiBTxKM1t3PSpqkI5XOdrBPQds/1ft4hLiI3W6GzD16XgsWPVAaG6uU
9fr4XCcK99namQb2Xwq88mXYsvOYM8rs9pYkv860idNJRt+RqoOwAgdsZnQ57ft6d1wTn8Og77cx
C87ONfT9UT1JnsVr+7iIqgTJXSZpy6XCVYRMw+D2zm5pMA/T9OKAkoaTB/XuDqLfLbgk0pH5icB6
AOfH91gHRCmrVod64SlDFRmgB+qzVU+2aG3FEXr3ct9JvdYFUuycAUSbOkiPyeA5gzsXtjdtjUIW
GatcmL7evPK6AmzdPGbe2ElRWwEOLkjVfPO8eI0eUE0h5zyVO3cp3oITJs6myh/4sPHROkvyMLux
RtZ+ElWZ3RuBbpIIG5x0W7ci9dcAf1HrDfPT+lCBQPgQ1OqqNW6iq2uAVj1+3vvELBDzKKWvZ86Q
KCHUZGnF51aGKmrWDqgqiurKWZwna7VkFteQSw0ldPyLj4kqpU75gMYUPLc6nZHFZasILDSxzmHw
zNJ3K6LiEPuv59gGja8ld1WW9z3v5azRFpS36vqNcmLhS0xkJVz0m/TAUjDprx/vzP5NGouJB6e8
4sxv1eWVQRa+vIRnuJew3M5juYs+688wjd97/0uj7KiwuNVmFyDgNHm9dimiDG7t2rOgQiA/BuFg
TYfWCn8tIEt4TgrdImAUmKkZ1duSgecpbYd/hlH8HT8a4+rojNW5CVrbIXIxzDs1YCNtBGoZVXY7
yiV0vV8MXTyw0hIdsQisJrrtQACPdeRSXVW8/zY8oPKOELkXU4luY9wtwJhep9IYbQ5PwwAPZNy3
jwT3TCvtyckjwmpNoqJKkCkgjZ7gootro9yetyBtGC5vL4ElR4uBAcse/yU0llFu9XcuH8vKHMWq
TxGwUCow7UBax60Ef4gx5TS/3BX4062tAH0VO3/kKdIDe1mcwPU5jWfviMO8+ml13LFTWGOzJH4g
xp9QV2SQB/XQTvP5nYWiW8TEzfIvRKVriCPiODCialR4ZuRpoyvXtYOaqd0MIqrlOiFTWbGyGnhU
JYgbJ8uoX1y506b3AvOUwzWH3m41/C3V/Wm0lXCQEIEyT6qoZNar4PlWv69yvnZ7M9jS+/atSgQ8
sHjntDve+cHGsv5qbdFZMZQIlJyqpMiAHbGD2jU7fgleTDFBLyJnx+lymDFjH6lDCnXnc1Ne/p+X
PCP6RyHHDlKY0vz5TYkOlnIcT7tLx2M/jnmVcNVJUJW0Qjz2b9HPmk6yd67haH2nBwBl7AAmQ9OC
0CpDJRxJI+4RfVs21wG5rHDxPGjqQXBHxJfT1IOymR60qqxcYJUcRTtubWZhuYbnhiQJhiSSWE2e
jgJShXHyQ2e9fmZxGTllB3TB7aLb5tSSfWmPViZyvvWCES8ZYctaY4QusyzoMHZoLcTbd8DiMPth
FhkJxeqTYgiNoDryMGq6UivUP7epiIeQgrlEDUYrbEDuTKBM8LdC5jQyTxMN0I5CNApxRf+2St7S
5XCoSYLAFMHj/O+mMd2xAWf7KfY3wOmoNEhsgNAzEWvDJK0fn/a721hrPaWBqB8ifsyG7IqO5kY6
8lBRvs9vDUwDFML38COErTFouPdjhYFC4pbBNrG+H3oUHAXb9r29CuQxeYPB1+bPHxObQv8ChLZc
hQS/w2juGJzfGLVOvKZ9OeUXvboRKfUxhHqLbUuZE8nn3AXAkToJfiFbfmOpLXjbzGqzX1IFMa5C
MkOCgbeV5LorSLqFJEYT3acTa+7cmwS6i9kr1OahZi051MIViimMN32YFiTmZQ2nWvbQlSmaZW0O
dQ1J4rNd1u/p7xedwG0AROUs5x2G6dayGP96vonpxLuh8VKVFJ3qfg+wH+Z4VRXqDqosy24JvD89
5jQJVVFI6Jw9ky+B2YZcY4EcoH48WanLroOmDecjMpCiAjjd5MmS5pTX1x/wRHO0UHZTPJwCvpr0
iS9hh7/1iGgo/rsycXkfO6X+177dloSlxRZISrldI5uAjPMaFVQqOZh0E12PCYN7QpG8XmQMojKE
nWN9eH7eLbGrsBGk7RVt+Grpx8KTpYVhvny+Z3KgUO+jZGtdWdCujvz+f+1cAe1JgJy1jnxPkXB3
00HL5BnFhHYrCh3PZeaK9J8H02WyLym2bQ+wjd67tcuedGybNeXcc/GhB36lIWoDwBgfkEk60f67
s1Oa1p6dyOhrEvProsalQYHFuMHejwJMdTYjTUhHS+IyycEaZHyDfAGX6qm7eA1mq+C81Qiz5nsm
7dEY+yIZ5wzDHL7Dgsm1ut1zdOTFLH464hKEpQL19Zq18P92Nm2L4jpt8BHW84kIu3MlXcWrH1I5
H/1SkrllnGmLoYO8bNdu7H9kR5DV4/culIZfERYUPqPi9Qn6BgpjoJzqLSk542PMVnACR1/OafvQ
hbORGh3eKvJgVStGEiUiAVyVsChH71gwRikmXKTcDs7F8I/nAT9BxFrjMVNXYALvcSYUVw+8kCFi
I8QeAu4o/gJ3gkHY8BNlAuwEUzCd+JyqR8tw4fKYUTjpRclQF87o3W4Ux+U/UdOdcOhflQU0Mk5f
bwZHHHqDJue03JSwJymJNw4/JikoKjyb/O9CiBedNwwSd9fz9xd/WSALzNJmcfpllVtd66GkhGHw
JxcJ1Z36x8Sh9JDeOl/NdMl2jC4oO5mLW0voLUbPA5AfIZccAQDWwNHOBjp8tnFFEW5n96l8S3ZN
7PNRvxuWSuuezhx3EFo1hyQfFj7GdaL9q/C7jL4/qxivFSomU8Ai+3r+65AyEPwmSqDyZiAc/oly
xppLZJmPcs+lttbbq7UUuf4IwQhcSR5hcIKRRFnTPyTUAjRh1Ix3skbq1T/edpwgI1a3+IDGksF4
P4Jun8+15Jd8H4fnKgQhrbNpTK7Hw4e5axM4/pufl5nvKF0P8J25bT98U1osoGmg4zgDZCeQEp/1
RjVWEzdECd97Af8j32ThdE4x+RK9hUPJncKTBOoFRJvWq5cqftwTlpO018IJOaGVEdYgSdlMJtp3
hPc+4k+0dnhMAdJYPa//Fbst4Naa/cayLjzqt6TeC2YStE157WpFyoROonFF393KnfdJGFJ1lcPy
TBWnLwDfGhsjC+yi8pbaXxjfXUWagC9kEjMzk2kI12T4mEjEbOJ/A5HPcy6k9BAlUxZ2JULf7DP2
utaYAa0iuTm9c/snYb/NH4zRbpVIEQINmKERFVG/arPb81CM1RfdAxQboaO0eTPfQPBR/O1QtQ1T
QZEtkK3m/NcFpWwJj1D5zkhNE3ePOnm/StQJHsKeilL2ZCHaQqWbP7ky2FDgmvT0QzL+nWG6RYdv
rLi9P3++CDwqzg5QrCj3gobEygGDLCaAm7nFDJACVzmSjFVYYgoRDMvip8Ynhd9zmYX4KA70HsxK
NLd4QAGJ6TI48eJ7EIOAVM13VtResOogw3kgVmcE2ntLrVHnfstEE4HnTtEUSXx0kwEeNquBmX+x
wtdSgzat8JL1d+BtpMSk/ps86PpJ9Q1ppQiO/m/6SgRja4+IMjiUQbKa3v1OBiH870I/cXGgci/g
624TGgpEXEWzDWEKQg/xi/jPIjddrzyHEsFnsKrLWrbj1iNVo5KfFY4AKGfV2htgH4AhQDPxoOVR
zgTyi7wmhS8zBXxQz0ZQCpPycq3hC5s9qWuuM9LzN/0uGpVb0lF4issSX+RxnzGSInofm6Es7pGJ
2M2HJ3tHPKMVFGdxqcaInNGrrYJoWATmfz5lSiWBwnHXL8AA+ryjz0PlG0OQu/vPRREHFj2mIH4p
MLu/eCXi0Xlgp6M/pMnPbfgg/qSAm609W4xndexnBJ1ejkeE9y6Or5sXN/IfdY/Vb+VojHUDcIYk
Y/n9eVk5DyPHHnAUahAttHSSNyeOqUnKCjh9aU3EIML5+PNm0iDT8kJ0uxxHx9BsEw2VrLb0cK9I
2fC4UhcQ76KDUVt1bDEIEBIih2M/j/VTpNR8LzplCDZdul5XUooLlu1vJ1YJc0UpYeQYjM4hUdGC
yaJsH4O5SFSo9a9AlyYmU1luxHywHUOkmuJkBggumIDXMccMgh0m/q8kBZOeYVl+GiVK1e5P63IU
0AY9qINmPr2tTxifWTsrgGwtFXB+MZatjEb93DKfny1bRzgsL5ov3qaDk/sq9+5ykxLhOFIRjcN4
flZuB0v7z5eoaPYcjlttMyC7eYJHR05Jf8hd8F3d/uwmXQP7j1a274Yb5JBwnK+DU+rKj9vB3v4n
l9EW5ymempazfztY7FjYGxFN37C5Sr7q3WzsCrcWkyaclCPC/LulqcyRXA3lIerzt/g/pV9gv/DA
2ov9rFpmXvK2De9ORVGczvrNfUA3YTUPjjgUQgfEcgTzVgTg/FaZVxquWUvatG0ESCFMd+iNg600
GOIlojhChG9yDnxmI4h5Khj53s9jvyUAqqTFAqFYPaae7pN2XqiXgFrOss6locdYj55DD048GU64
VF59T1p5Nzg6ANGgHUKZ3p9W9iErGodxJiTY1VOWORy0l4ipmc9J5l1Z8Qq53z5RclQlw7/BkHig
63HB2A0D/TeNV8TzWWlgwowqNlh+dUwDHdlzHq1WmxRJJ6ekAPceI8j3H9AgSI0ghiSUqGJhk10d
+nxqrjiDzNwVd6zq1VkTTNKHlPqP1b/hWUMYHmHvADi+XQVYVXn+cdv6NqF2N+YYhJEO5vk9LJn0
Z4dCWSDAVriPV9/atOJ3G7Ldnl0zsuKBIgbIsUIVj4fdTMC3mmX/qfpA1wQm83LgrXw778fF+Vpf
J5aJTZCOvrNrlSBWt709HDEtU+1ljpCeAHozn8hzsGR7fKwdXMa0u0rHiphUdGFWcOoMPliR/W3N
LdyXjZoq8c/lcXCV/WGP+F9x2uV6b4/owc3yTzbFwJj8dADKmkhhNeLVve8+okZB22cOQ6Jdca8H
Plf4uudcZvvYmA+ZAdu0HRO36ZeGvaaJI0VG2Se6zDQBKTLfcXYbEFIijdOE092OfEgtUxiOcZvV
rop/AFUXTw1Vc2KOaZQVN4OMeDSgMp2WggPutYtvWWWhRM87petX4rqJtuBnRQYz3lStiaQ196oR
z4MuCnPaVtSU/zEBZLDFM9yO9tpalz2q7WPHS4QKJUM9zKl1JMz3iH0K7r1oGZAWRTTuWGu7HjVA
V7SKG0F35rSisOaISa/zp+HGwOrW2RjasbpYi/1/OuSCtXmOCS991CW2caTXrd7GPgI9rDFNvNkJ
DAGVTONFezR652Vo8OaeF95qWW6vVVMLUksq5p68EVEBjBaQ6mxeYriylMaG9WEDfmWlY2+myPSA
qtvc+MmEwG/0BwkWI9PwBjOCe7ctfIdyYqbq7fNlPLGsEP/Z6xJpFtlUBk+Js7eoDBVlH1JjNbsm
f09mpdi2kfPT93H0wcJYdUMByRwoJ3kKy+txfNJOnw5XreKAViiAi5DeD4HPkac7yjQUjvi+gz58
Z57QUSYlclehvO0lVtrEMqfEukIJvz1gdU1FqjLPogC/hF6cl+cBn9rDGRoQO9okXwUymIhf4Ub6
caj/OyKXhKVWhOAPYyRJYn5+pBzMpKxhdBWQffl/H1jd1llRCxtvLVEVD7sPBIDqZJofv99L8+sn
3/+ol8ybXd8i0TRvBfAHVDLPrJE3xFiPpL7Fp8geNqbRNvDkaTuNxiMScFaCkrb8mUF+IRzVaO1W
UFLtwq63NGM3FJnfdQBpzyMFVumbjuwhg/8Jjt63M20qN7jKNHOKx7MANgisqPSE/ZCYyYtKIOU2
35R8+lIo8jh+GdVH5Z4JzUS9gGtRoRED8U0NyPKIAMxoJc284w5tQ70eCx4TsxMDSt2AjnQ8pdPr
sQtxg50bOKSddcANXM6pVfDVTUJTygjo0JRr/CPb1REYuYR+qbEei7RrghYB+AfIbl5981hMzE9J
hnBdUbGz7pBh24EAzQHLhNcB8si5q4XG11j0Km5+AdD6+Pgj1+JkhGCqFwkckgraVWpfq5U/E5FU
8WM5B592yvD/gh7Pa/YfdPAfMshpiSiIrLuN4DVIhvEtWx5N5zlnr06RLbZr9Sp5F8/Q/Q6Gegow
D4LkI8zdYnVGUESvApasY5DN/1e/Tr9BBiJepjzALQfVkLOGn24NE8tWeUvxk/hcpaAQDh0KH61m
j/W0LTulEhQhLI42cJaENodVoby1q81jFDLuwwlMHz4bun+EoiJDhawd/hcDmAIRgWYQq51j06bn
UWY0ENlWXLWxX6dfOcwjuu6tAGqzByfBdEA1UkEs/rJYfKHpJJnJ8xj5p31ApUogRQ5G4+rxeZNP
ruCA2ww1EyPLq3kQdx3BBqQB900jt3X4jqrJ/Sh/QPNaNNwnyQ/+3kBct3TPDPO6WVReFo6+FlJa
kE7I2/u1fUxX3Jd/5293p4B1bHOL6WwwAYmWl2sck2xiwXJJrDt2cMhdc+UPT9yg8D/1kRHcqcdy
vLthILxOnnCRYkqhjjISeh2QggRydWBp6jy5WTqty34qu681PS2phM/qHgcxYfkG+qyKpho9gUvv
2wU0q/n5IqU8qobugaPB9EqgONyZ8aI8lS4cF8FpETTVOtqVShAOADiN5uCswW6LXN9PSNp8ddCT
AXPcO6btAwmnyLwybJe8Lx9GLCPPX7Zqd1i/MC7zq1iCCduvFw8iUzozk6EVhj/QjQ3/qMw5neT8
FfuYmPQw/N9tQryEZeyKcnQMiKjrwAd/SH/3OdehYWTgy0yekHGab3t88g2KUN01qCEu90cUvnkS
9su5CmM6jQ1FUiop9ackRYmc+fiyXbEs5duLj8pYdbxKWFLJjA4soTPFtUibz54hI0jxMMIUDrQR
dfswAWWAogoEhyrjj6GSM8FUeIMgK2GkVpcm16t5JOdLzBAPprhxVKJdHJJlfdBH89j1hbcDL4kk
OW9QVmidyo4sZ5JJ3JVMPi3c/8FCuFb1aApRaEZsLDfJO+q8x9NKf3WIyvkM86XW0rVdr66EfIF4
ghmhlHhzdkFgYNeHD9y/i0dsNHzEHmRJz31Z0BNYXN6u7k3It+NJE8JwcYqMS7M5xVCEHLiG5UaH
odZJiawALqM8mfa+XWnXLm2dMN8H4vOiFMTwX9BwYk+bsElaoVenilPUodLNn3HcuYSP4BZbW7Q5
57YADS8YUGSI9GtXV4V0RRL24M1g2x+PSwwSxrPJPw0BPbGjyP2IimaPDbzxoxypPS83V2x8Logd
188YhWfUcNL6r12mbY09yW59+OLSRaPbEzKHJ4QbGCuvO0MvxA3wJAphAH1Wri/BiE6BUawW/kXG
Vy+6WrDpbJMGwO2eBru9UiiNviliNv+gpQAWYaVL+gryjn5OF4/+kkFDBBKYL5bMDZOFRno9fPE+
OhQ8nSZCv38s2bX7ZdfmCm6NqNpzRCgyjl3YhOa8rsYuLK6NtkqlE8f0wqUnYwehMmkSLRqifvmT
HjFItMXcCVXnWWwL8/QyAyZazq9sc6i+hMmK89krbBvYCSBCAqH7jHMzxCzk93OCNkmKNAcQp5OY
91VFq05g8PxUeK6z8db2KlLd0+CRm8qyVrrm6fpnkoyPDu+HLTj16DhwGueoMistANksEQgSdHJo
PDsklNSe3p99tk1ROzYc0AAsfFnqRcRUPcuuFWcP78nfRse+zXRo0eaalbEFFovutPyUAFZ38Ch8
y4SSL5T+7uRb9fula+9vKExOjyxN/ClmDXDhK8DfXR/aHzeSHgJlUX/O4LyleASnDz67ydsmvLIC
z6ftZLPRqEJ7CbCYiY0XogfRaFfbifWvyFotT20ezwOQKmXTIVeNnGEbx136N+GG/1aUDe2R5Y71
vONRyZ9dGbZeBBa8H6aLkaIxWU6EhKJy3giB+oVKZgOSQSb4MNEtV6zNqy8WQD/0YBc+9kce7VmC
soHs2X1A/UIuDiccsWbrKev5n5RFc1yWUmXkzwshrYD/5b16aVr/dKWhUXxU4ZsBfI6dc7a5DDnm
dVizJr6t+G1PfoPs2fL/rT7KYDFo0/bJjUDiATJO8Pb7w2eVX477sJR9UR+h06ZdViTWVCa9As2f
6EKzjcrcR9FEmlYZdv4XOXMnLIkQcr+tZFATg/4krmJLG4rqZxzQoz2es7jrtTuxZj5QTeoXOMVR
yAQnxt1JEPdxATAChz6EYtLZBTo16fo5RXF5sxB8Yu5DOhd/XzrtHwJkxNMZ6d1KFD9V70X9omKo
GbAPT83uKVWIBq44f4Sy0tdfX7SYYHjFAlE3pJxp4bEQ6HtGC6Zg/KajC91C/UjgZAoFi1OX7DTG
vrcfUIu3EAwXo4cqTMOuPRMS3TQQih0kBVQQryNTa2Mj6r4fKaMG0FN4HunTsGipbZVEJrRFBRha
5gTUCiClZR6S26TG6wWmfkRxhn1/l2sYLsyhkr8/EeCMqJKMtO7fJR39oqAmsoDh14QQwqXlZeNn
92GpuJiO+eRpsLd7JS+P1/JWJZjlznC/clK1q9FtkLWmDGqJ721WFMi4TnY6sc+CsKZ8xXIPZN0m
EdWKsh5wVyPU2aRkgQKlXVm0j9oiRIuG1/hAsHiydUlfHufsDEtjoeYUhSYLo7A6C541aBXA/d90
4vssf2Ja/Ma6HiS+ROV96JVLCcPu7VbJJGiXbKvC5LHxOMLVg7ea3yTrkpThREybzQZpsuUkggb3
XB+Wh4zUGalrqPmHFaty+vKYDIQtG2GXhvop8lIGsdoQpAxv8gc+DlM0mPwDi0J+fml93miR1VHl
mkV20Y5tElTx565GpjX5c87Nl6enQdgw0jSpmy6zAp7v+pO4HjzAeo3vBcqkrkctvcPg/ZL04GGO
tzuI/iNxHfcJDswGh9+XxSxGa4c2gTSIlWkLL2ruQ4o144U6ujSotlZ8ajAJVX/4ew+1HuWtAY/r
t6N2A9koXXnaTtNhMdetF5cIuQZ0CEhvzmdHpsrZNjI1AD02q0MNEl4oypqilfqHeoiVYE/utkjB
3OeTniMEiOOWmc0jV4ukQDD3Fe1KPf7eHCyr/X54gpVZ0YyYZORu5y24jD+L9wtHWdjtMDfzkJe9
aMPef+nvJ/j3gFERD83W7jT8h288KTOGDWiyFfh4/i/AdMJMNTNjNoBHSPR7Hmt8F36ALkrdefXf
dmd+iSaLNn5Keaa0KRmJKQWqy84oiOxkKCcot+s4BTe1k4OEkFalS9DKnFC2bzD3WFFhUghbqOH7
+OicX7BX56vXfMzqPRd+1DZiM5+QP/6k9EWjuZfY5dwpAZthY9bnG9kBaUPNbqguQTpiIXGztSIw
Prrrs8xnysr+iIRpTlmmJUpnGavDq1BzkDwIND0M6nl7qErkJRlytpxfgqNzlc2/A5HwDW5vTm0s
ZCzsJO9cU8s7KiPXcHHVcW9S5SQuHNfD26iD2jMyqbbnExCZZPIexO6akwyORIT9FWXC8miJRRMc
O0XFVRAEAFH0d9LV+Jjxqs5o47yN2dxZ9NwLTn2uyOvPbAQdXL7WnLdZXBkp8Ug+wfZ+UCnwcJuZ
qwRMgjAJyObL7NCbUaXARxf/B6ERzYHkj2rM27ttmumcZ304alN9XmIqZsY9WDxq4WkOzmhBJrbo
xPZN0XAlEqHi7//a0aKq2W7cCzr3uLyDPhW9t0We/F9r4pJ2u4K3fMtf2ZoeLfy8yixYvqj559+e
C5Osb5OPvDcRPooMPZ5UhIG2xZayZfTdt34Q9H9m5OqX/OqKW805PgVN/SXzeCOwWcZO6B86ebBf
tZS52CB6fqTFRSg70JHUgpASY5qfHnjgZV7cfk7pLzvD2Q5Xxkmkk3JmXzjBlNW6zcGuXYcAor82
DkQf2F6VvtcvK/7Z/5nT6VF2rj6tFHCVH04RKSYehvvE2vnT2pS+FE090x0qZQ9/Q+2xieCpCXjO
52yEHbbIjMPGCPqpNvwKCauFZFpPhF3yFrPMCcewny+STo1LsaRt3zliCqjV6Dl13gyFecG52E0z
A8yQdM908a0dzlo6A/tGe27VC6gyGlJmzzzyyxAERgBb+ER/df8BOM+8pWwi1k886Jy/tRJsvfqi
wvrtXyIFPZlutbnCz1LU8E5+4MPCtDirqUijLF5CoQJ22rkZfyWg9WP+4RQn8cRCt4O7JsQDlZYh
sYO94fRo7nAm5c/G2zJOYECoOl8Eoanp+HNCICB6vfw+M17t6KBwt1NYHCkqg5Ausy/TFic3yjkZ
gBTemzhgo+1TFMOlKNpGVKi8kUJLJFZRo1dL8D9fffGolnIHwIE2zmateiDMnXbQuX2PjsvvK/U3
gfcODBEtgVezVUDALV7kRbYDZCIPYUoK6MBnwaBk6ECPE50i9lSPQrzpsKaRB9XyyQHihZsUusQj
tieNFtGAUG0cYTCclYGtvYhVIKKdXXGXE3VJ17neNsELjH9YfgRhkrFOQAdeBZI78IBXptm0pHzD
oOUkA1O6Q8vNBi4CbV+oNigeFwnuJPhit4m6Ch1c5OAHZgTN+4UnQlkuwGvsjF2HnjYE55MzzRtA
0uSiuKlGYbxB+0XYU3BjADCI8Qo9tfQGlwxZBegmCp+z41Qh6f70oJhkz5/Sxs5i0LzA4cykJ00R
khpv3EXg8po9I5+95T4DsjtL9tm7Ul8RW8u3vXKDdwUgyguqN8fRus2a74lbwuEumbAfj64qY7w4
LiHkw+DCK02mGvMfFLS0v9N7ioLeBxoM6ade7pdY35Mq1P6s0ATeFY8XOysMgJHMFsP4ikUQbnvd
nurPg9HqpQdwfv7V88GDcSntJ9lkp6U24z0VszYFXdrQbZoCKiHgbDIL25qdq9lIeIromNyYNgG/
5ka+GF8KonjLS22aH6R0jzOtg2OVatxFmRcCl+IsVKrvcdtYxzQVk0aJs9SWv//9o2aPXZJESBk0
yfJnhIcdUjafFqfWiMr3K7cM/rK97vjUXo0qFxXZJOpx1KSRMGfVHjktf8x/01XCo7lgrdpHd44M
4OCFr2LUlkWyXc6xbNFztVgBtE+gx2V4ws5dxAvFaatxKk6yPfQuioyi1zubC5+k7vFiqHaEf/nk
4ffitEgEBwwRzfiCbOo2LCuy6rHgEEQLvTfi9VL2tSH4mS+E6rFcnxFbCNu27QV5pwCvCAraT9eT
q8WZtdYscrHFb0fvoyvKvgMKB6EOeUsoibZc/On5UxGeg3nh/rr7OlKFHZUPl3NGPvO/fPdA9yQE
OcCXriW1nhBT4CZuP/1dPDQz7eQ4f2RWxystHld0uDhY2pb6XUwC+JY9RG7ehy8/xDTaxT4J+Ikz
BfaV+jzvUVMe72BqNibNC1xfkycKjyOBaUai1xbNWXZ9dldXZII4h/+Z/aASOSn0dpVKfePMmPdr
W2t1fRzd7UoSO32Pb8zASfRNZTLN2JaeKlS+9BiBnvQ/tihk8yvpHnjehiX2qcmygFH7wL4JNQJL
j6ba1/wXa4vakcUg/xAlOSH7urtZV5auEjbOsaL1KYJ7sLaeunJjB01mdeG8bgO5TGPWSujWfYT+
UZsMtkhLhA14U9FYGqtv/7geeZZzWGgAzcAHTS0XXIpMVBAH5SZwzm9TopP9CVV0uqzR6VsuDdQB
srw72TVDOYtqbt1eBtLcg+9RTpMqLabftQK8MvXiP7NPN3A9S1+mjCSWyzkA+dHE8jnYRkq0Km8z
QZOYghWjXOAtsNsj5Yt5ZyM71fx8y1hFs/DIIRx9/QvCDg6F7GUjQSIEuBq6LSltljAFuMwybnd5
SmYWkA9U12aVYf2ZS8K7pp/nlciWAuPn183AvWP0GF7kal2QvIzwYkfq3aXKFKJfKtAmjbXDuDKW
lJYAYiBY7kDzF2n7+W/zvpJibNe2VA3syjxJj8KhH0iwTPRvwya1s146wNhH3EfZFV5gxKYqLFUD
9YIIcujI/V5Oe/XeT7PH4tAsYosVevPUKomwEqpGCgA29594AGCbEIYZlku5ofFueke6AN/2osJw
YgbC25nBkBAMRz6WQn1S1MZhUoF9JAyUYJL3AHBMtg9ZYTgjb132WjVvlpU7rZXMRegmGl4ELkZB
rhkqA0bSVZ9IGvENdo2F9JbgJWH2/wGY/avOc3ud5NIFTet47s/XUKahqYEwsTL+Bplg848+EFSc
3EooOVnMS0yilFfAWiOaqu6ff0vSBeCv0e3QeT9oUHSJqZdV/k9FE6/Rq/PLRG/wHMZHowEW8q1x
gI9D31OwzI3oOoZmn0GVj+SaCQmfRWBfqsI1fwgRbAK7WT5eAheu26+w6/HzmKnmkHgcT4YPvQzQ
G/MT0aWcCtaZDoRD5UqQGxXPE1sJcwXd1ndS51F/uxLOLozH1kmcKFwXHiHR/qWwK9leB3xeF8FK
oeuxeQqqGYU3Ktq48z2TgV3RZDn8jwxmffnx9Y2SXHR2Bx9qxH38EK1cQnK71jHccI0Ed1cT6khs
I6UyQSRrZ+64/+wshLwmbFURfAf5rXgF0NHv2D0P6irdSOeDt/hE+t42QNHsbetueV4oE3cCsD4B
LXcofXbq6+MNHnAlDdtD8SnoZYNLVtLlENnXN4ryOk4MbiAMK4mFrMl/JQ0EzV95kl3Ozmnz/WO4
0n8JUDgR7vNKMXx0gA7Wm+lZiA8tD3fIJ1lkEHcQHM40jsemE65HQK7+H/sRwUin3yfXEsUWH01J
skJuDCZGRlnGQ7xjWUrO7zrnjEMjFT+bJMGZWauWHrFFTkNEB08AGVi3qF9WU1DchqVJWrDVVlY2
CRkmooE+2Lb4Mc0r7LRDLP2xF3S8fYbZ73qPLyubH2PwnYy8xIU+oel9iVUWv3pyve3Wl7+w022W
n90Yxb7heOOfakQ/eeiZ3AFxZDcsv1B8/CWr4jy4eCsIkU3buHIulO+S4Zmqmmhm/zoFOBswOV4F
izmYsJImeJANSvu8OgrTSRjKj2oXO0wVL9afUFQ04dzUUa5ykTU/RBbSjLBxGDSCyquh/rubEdws
bbdhUnMGKHaAx2wpzIR5R/tc5QydTS1akqT9mta7mNNzODgvkiGulREdpsk/kwhBq0yvkkQct5WS
U3OTYC/ZaEJyb4fO8Qextuxm9WGJUQPaSuydMpXrhzUruPgIEtASxKEWpl47grtfHg6Ff/jzFHaT
831mBG43RIMjCyBB66FIlbXqqagLAumyjqpt8sDeFLHJmSqjV3slq7EgEpsENO4UWLQsPzLjKEHV
Nui1HtxsO0q6jdPBn3lOs8XhDloD9cmaWEaAGWVNzj67QaRw9DGAJ0Kjk5Isz5EK2WQBAMRdwanh
DmeFXZSD1FO9HgfX1nI7PdwKhZLZc/IMMDVJ/LaqFld0MvRmpQeWYJHalV53KJIvSksaWtCj58fs
GeyaX/YBD5I4sKX0ioHJEOf/diXmGfQIgsxKEEj41lE2AF5CZ88PRm1z7O6d8Vwmxfu/kNkWobaZ
81mR0qDKXRhFvBaSmSeIHZTU5kh266Dw5z/nwudoLdC4L5TsbqlnuumWM0tKLyIFa2QQ7WUrD5tY
j6ppzAL4wcWkUgv+9zIsCyEAyI2CJnTS9+uqpRfdPNW18klMwo6TJy7T191FBmlRzBlLdkJJurnm
5NsBi/hzYErmCOJiLd7PbmcTQswkG6NpXrWcUGra+bv9gjZ96HuWxVuASqArjwDOxtF/0uy1NqMj
PpaFxWnyr+UKOqZYcnZrIocn9BuHskGDIKSJFg/LK2ZTki0SFkbRmmbf+XD/vMA903dyidCQIc7S
qywyU9vQMl35erAQjO1BOyFBs4c62BASh19SQ7kYYzO6MzjSkdRy2EDeAVAQ7Aqsj/LdPLzV258A
etbGWGwsqKzeY7gWAdBtsFLgG9vRoKd/hZBc1rWWA6uHxpKelgkkRMMaVxMf04bqVE9uD6KYuA99
7tQevqyi7JGOUIilSnTL4AISYYkhOerchjXEKcgZ8RLlCr/jd8WiIgtFTSYIbZiUYboxO9K4zUaE
mBKyV7tup0aR+a7Uqh4foho/tu3bx+AGvRrFEQq1npFnechrJDT6Oa6E+MmDeTyN79oEvZk9GGdF
+gqJZUXVHtMOsRq9RX+P1LXk/2s0u/Loa4P3511OaY+xe98Z11Kikjg7lXXYoxYAoAokr34NC68M
86AOPxWUD/OA8h0Hw38bt2h6pIgWyE38Q550LScyBAsrOiXzMzthrq5P5aWNZZhmil8hkrUTMtoa
9VLp1zufPQil/HSOLYe+SLjFZM70PKI5iUfGR0S4qJiODFAPA3jaWgdO3Jz5UnBWNcoQ5hNc5ROc
yMKQ0DPqCBLaBg3rL1ckK9fyKnrwP6QIGTpI/2t/p4mCL22z8gTkAOGzdEB3Ylb8dxXBASFNpqJ5
+VP9OSZiaA+tTEi9ftaeUK6Mho/I1bnyBCmrOHCTUwfMwHqHSr3Vx3oDa0ecTS967rt74lbk+5LP
7wJiqrDCvheFQd5yr9YNPyuHz4T9WRTjn253OsHoEx5k5wF4XmUxGwUI4zyRGb57rNeOkrZCNf4T
UGv7IWw/ZNLNVJLItX7HIPRiOzCGrHh5Dultk0/DGV6lLdT45wrtFprlXoWrz7pl88BKIV6MVHi+
0DNHgXeijuGear8TI69T+vBbMfdV51Bqezp1lx004PU5WPHo79j1IH0RspXq7doW7CFmgxOPRd4J
S/UvwwXUteVXIVwwzgZjrbWtkcPfWy/I4S6HY949haiGPZjGX9v4+6vwKtyQI0fq8yOKoU3ggfM7
u+5k49Y7QvkSHpnLRsmciznwGtn4qll6dyZOEbrdqMErhQ6gyGg5b9Z9bhENL5PWh/5U2nrKvYSv
XJIV7UccDGwQi00J8xmO15t/0wYTUq/HDmzWYMD2GwjVxQDzYxSX9kz02WYa9pS+qXWnGZOnZmoP
5bSAPjNu/iqkqfnxViBRN4uWDtRCO4HiiiXdEZzD4ekEVgYzJ4RKdk2aS5JukuC1s0PJeXaJOaE6
S9DO+lSIeR/HTQNLpRSO5DVtt0K283Xg5yr7+TKouIxUvAkZ4sQnU6A1sL7PCHkAlRVUGeRcM87e
TIN8REYDI4vJ7F0LKb8W2dX0RY3hcAEpZB+4KCH6bpXZv/v3zr8BLx0v+wFqUa25n3UHy/SBdGxy
INgi9isVtpozYvqlgyMTFFicsyoP9jE7/6X8Butw1CcD2v54PPDARpryaLCqWWUEp1M1xxlpUTKl
TBcx7vVWL4T3wzm8hJDh+nSZY5M4RWFx5TvGs9S36jF4CytRrwkc+O84G1jb9ImL3Tv7z6T5FRrp
0ukfqRZ223T8RMo0xPPczBkVBcfb1Zkdls+cdfMS3mWYf0tHnEfUQ9g2ca7OhZZps+jKC+L5BJzd
T2rttmxCB4gwIGR6v4FTMcyxwdTzg4ZhRYOWft04L+q2BzGTzb4TVEY1h88Wwm3G8xmVe6QgqZCe
vQGsng1L0XyyZBk7u9qGi3Ndomn7XOSmHG6bIIyZVoP2bAfOVcXHhlVxICs5CXYzN1me1vu1xuEg
D1SDCOTNYGgyAwRkR25kICSCTL2ySJVmlRAHT4P9QstTmfZLJvsHZxWTHpz5gM8Q/ghFBswInP2b
oFKxyhIGlEJNS8XwHYP3E/Cb1ECSmd6AaTyz8r+pNZMr+sPL2quCZxuBZHi6GpEPZdSqb24KRGcW
mJXhaZGMhfcA6XXATLa/z3UBwny5l6/p3WX9E9ysxcru8Yyoc1YQ0yIuS7azgwjcO3khL7sVCFR8
wQrmA+5Q9RKPgaLon0Ln1DfB5DTsgeHo1uuZ+axE+8u69rUGaMxcAJXC7WpgNuXpOzY5e6ELBXuR
50AjWZCVtgu1+u/vqpE4hmyewltVZ3CytSmNPHPpKryDwdoLkTYXddWRWtEHYacVF06MZUjHg8rE
4uhJMko52azGlfdZ7m9TWUvfElXyxdVm18EaWs5ghGBdL4WC6VI4dWIeIpP0/3e8QPY+H/vS91Re
t6iYaR06/4JIbDKTARjyubsXTgqpfDD1GHRuldmlormq7+ODd9tkVOzXi+P7oK9xCP1myQX7aUE3
gw4PM+ydkKZfYtL9m4li1ogPPyw7tsuIUV4tVKFOnUcNwDypDjFTYI1jEwAATgZJ1PwwLBYG4AME
DIjreZ0GCrcA8kfJLu0HXXU/KXlj2RYp8hOnN2R7F83l5CKH0llEuqqwhSqGI82P7I2V2DN27ow7
wwNeXLRtISKiPJENUySRlGLkKd7BkWOYvjyTUoYaxNlEy17MA3BPsh/Jyy/Z8MeTXqut156k9mIg
gVcJXXPp4+hfKyre5isQ3AT7/bjpmkCveIGVtltkqsQgdnZZkoulbAIgiSgsQUOwldlrkmoLWPHt
mWPePZ1yrMmKxeMqJ5wtUj1+6IhUw02myQWSie+iVQaNJWerfbK1mp5oDJBv2EgMJXuoWV4Fvp8k
ur8HsB6eAU4fUXpSRnBX1XYR6ymfaqs8mHI4jJyAtbqaqnyT+rn35xC06CeOZqlQE4rsX8GAgmVN
cAN35k2tuUMYsen96RbXIUNx4u6MZnofrvzNecSrJI5UbJRUg2/gT6DhrIMTvtGvD1cJjDWX3MuH
N/KkiqlS3SBzKc2JkSU0EetaAnks1GWZhlxSM4ba9iEmOJnx442kSd3D8BZJs8/LIZvPsR58LvZZ
RE7233Qjqvkk3mMyR4/UI78Er2xuyAy9/rSYK+xKc+7SFK99RZp7SKGCYVAFAiwT4nGtvrBNRl8f
CdcbQRnxRnByvoLtQfLW2Dcd5oVq7SJZgvv4DoxGUKwGM859aZxyhZKhW73ZHdyk6A7YJJhRSYiz
Mtq1Olh3GMmbUquRug0NXGM3qelRwnaS3mArdYffqd5oIzza/fxNFA72WcJc4RmJjwpq13oXbKdk
NA6vztDmzOm8hwPgA9TZero0DXECtbI8P17lwCRKPdNGks22L1DKsRDLtUVUDEqWoBCuCh0MmRBf
lIt+qlji7QWa+mqsubXcNTo+DeG4vFNpfcmU3RuhXPCidqVTekycc/AMVu45BmzQMIWySRB4q+Tc
1WCR/+nhauHhI4Tn4wRQdVS4XbeXPihhQoifyQ+NerCpqh/lxYfYQJPMS410w04CbpLIMAi8BQ7e
WToW7+quYe0xLFSVerX7TpeOZkaBOeZY613vUmhkPnO7I2gQwdIOfH6ME9wIOMq7X5/vGKtwNJGw
dnaPo+CC8REU8ALwaFfB7SayFzu8AQ5ZRHkRHADLYNauSJDmS7w3LWQPF4beqVMbXTnrshg18iO7
SlC6IRmkpEKEvv+R11mw+N6MO1NWUEkaUNmYBJf2VMfd9/R4YhgiN39qJi57WwaFYgKTe0G6iwgw
PgxNu/tqyzGSonZm+M3YzXGBZPfkIEuaqeROvt7mb5AIReSX2pexKpQDVE/LAL3LEFe5coEZBiEI
tFC2p6zpB4N1uMzhPJTRcLw56Wmzp89yrIF8fujgSoAnehtiAQmBYPkgmoyeRwFHrx6b7fhqPZBi
vGsFhqqLZKmwFXeKB6NU1cCQosE1q+gROKPntsRM9MKk+KKYQ2Con8GbvgjM5DLBTFKyv0agFc14
y3mYbbXr3wj31/VzgceyWDavGnyFPU5vVGwtKjil7e2QmZttmuJfXgr/Pifi4pCQEpitIFgaTps3
/LXRc5BroIzAeKQujkU1tfYq5jdUNoAChjV1g76dy51pfpf+fY1kTvINPVEg1wtJ0u1wu+EOD5l/
CNnDRQZFoTtELxwhP4wzfHW/+dd2RduBKXjZyrgWKtDmW/o55OqjSYrI9+wgpeN14D3R7nuKwMMX
7QJTIGy2jdekGmB1HKIarkjtdVjqWsnaSFKL2/xq7RjnrTNNUMrnx+5XGgdM/l3/KCJS9SevB9Fo
vuxHyFPxIH3mzrHhXHbPDKNUaJaNqB7A59MdnGZ5Ce9pO/c4ZNveWrV38ymh3lFLTYyRoenHuDWG
M/VXRdpbGsI9yDR5Vfdwip6gP0+/tVCB2yoF2+9DDbjg3ba2E5CWLiFiqOc5B82ASsEJg5ZgtfxZ
dMPX2ecQmg68/b2pa25Fwcesm+bv9Sda2XJoh8RTIIEAZwIapHsaaGzzBqQq00GI7/UHTaLPa3fs
8EdORd8LlESTRSRDSaK6QAgjSKQ49YKwKOeKWc3Ep+0Nf7Awz/LkpXA/DdcW6DuyLF0Bgxv7hqbe
YWZe++RIvcsGjgxrRnuNoeOXazb+D+1WIijcJGQvd58JUSoepLiN6itVoLujsE8He83lvySfPcsF
+wDt2ob5jW0pKycrmkuKmI7qqFyItPO2AA5YPCYRqaWs4Le2xZ8x5bYq4ukbSqj6+CJk0MrEunkn
qOK3ENnkX+tSyHOaBmFs+yi9nLxbuziTghBcbdoSFZmFXsn6iYMRZTxxbbNbSOPnofTmYUsZp7hc
rQ3gvjGqrBKaAGuaLVzzCHbUDxWkhMXpUkUkjNVTnEOxaD+yryRCemsC1UwqbUuSdSxLuuvAK/wQ
3mNBxUo0PqVolTS1yn2PfIq2oiB9W96ocUl5rvBKPatTxWacELDM09unaD3FizPF1UoLOSuY2vqK
IFfeDMYvcUoYhaf6/GxMLfgBnrEiohDTV/3t6w5AuwiEJiSMp/B+CglNcuA+S3RpNGC7HkNLCOnN
h+SJJT8gjhCZAYyDtH67upea+LtClmGXKkONK5OQIE9d8AsSpHMygsEgCUOaHEIRpfh39T99qspA
FdTrwLjpnLz3MnUv4eMv2l/Cz5uscmZRUT0jbcLAyLonpzfHQXAVAaLvDH1Aar7dmMM/KbI6iyRS
fw3K8dH2hvQuq4/ciRh3EGnh9Chpl8knRsLCl4rrCwKYzC8//vJVB6mCHwbnP2TlihapbDmagobt
XxAcztOd0wWU8+pe9M4yZbyCG+ODxiWD2V0Eq+i/JJwKb+ovNsDq0qlpJ2bVECTspZiZWkNWPVgD
KOhjvoMl/tX4v8TMN0k152Dm8zZln//uWeA+eV0X6BAKY2M3Ed5QGhqrUgaAlrisS4OUuS1hLFXG
wOhQA6Jp0Kr4erbyyRYLs3soCQhQiF4Y5fJT716nzN8ZUmtmJzvQ+EMYmQUdsB4BLr4CcQ8Ra7ii
BbrMcHFg6RoxkZSbjs/8a8FbkymnuK/gqjb/Q+Sja5ckv1w4BIw0KGBO/55syidpVEYbB2Dq2Sly
r+LMI9kdUwB7xh/rrzPA3foPJcNC3x+wQIXXWR3MjlIxjB89tkc1m4DDpLUNk4XhgMxr/mPpn91S
r93G7M0Ta6EXNkkUfO51YYUJeXs86sPNtc07668AsVoRSf+WnPAW1nYOI1+pW7pKYJM5BHlLJZuw
XHtVZUAD0sccMFS97ef9xMznh6n95gcDE/fF6yvrNbDE0c9Hdo9AX0mNV0y42eiohttGSxWFoWVh
9SK0SgD3OQZ7VqY6dYtKvkuETvUyVC2UmTJiDm918C0vp8rZeCy/3sC9S5v2wE3lJlbUJjnrshXr
Sl7s6tsrIO3L+XOD6lyB1eia+FHPyDTWUzhcJzMzsa48Z+CtX6syVv6KYlgQ0SEClu/VFoCbh2QO
bpzuik3npgZu44bxkMsYtnWbZCBoOukvxe/F/UHKRGV+VfAReDcpFMhdybK5Dg4yjGb6yRhX2VjR
7Y5Q/Vsu2TaFkKnB37KFOpTsYzfgL66ObNoX+dZopccIGKsltzbuBJ4r4kL3F5BzWBFwxesuVmnY
Aph4nUpdyKJw9zfCf4oXHjhcV2zvP9OZelsqeel9dAc1XijVicPOJFCcyIC17xgwENX3FBY4IFux
m3nIpGexLiamIg7RE4ZzpF6ABi7DMK8Vh4Lcdez6R/F4pxB7537+mra34AY11V5qaDgNiLmrVw==
`protect end_protected
