--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/
-- ==============================================================
-- RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC
-- Version: 2013.4
-- Copyright (C) 2013 Xilinx Inc. All rights reserved.
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mul_zeta_12289_6145 is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    data_in_V : IN STD_LOGIC_VECTOR (13 downto 0);
    ap_return : OUT STD_LOGIC_VECTOR (14 downto 0) );
end;


architecture behav of mul_zeta_12289_6145 is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "mul_zeta_12289_6145,hls_ip_2013_4,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z045ffg900-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=pipeline,HLS_SYN_CLOCK=8.160000,HLS_SYN_LAT=4,HLS_SYN_TPT=1,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=0,HLS_SYN_LUT=0}";
    constant ap_true : BOOLEAN := true;
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv12_0 : STD_LOGIC_VECTOR (11 downto 0) := "000000000000";
    constant ap_const_lv13_0 : STD_LOGIC_VECTOR (12 downto 0) := "0000000000000";
    constant ap_const_lv4_0 : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    constant ap_const_lv6_0 : STD_LOGIC_VECTOR (5 downto 0) := "000000";
    constant ap_const_lv8_0 : STD_LOGIC_VECTOR (7 downto 0) := "00000000";
    constant ap_const_lv10_0 : STD_LOGIC_VECTOR (9 downto 0) := "0000000000";
    constant ap_const_lv14_0 : STD_LOGIC_VECTOR (13 downto 0) := "00000000000000";
    constant ap_const_lv32_1D : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011101";
    constant ap_const_lv32_2A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101010";
    constant ap_const_lv28_6001 : STD_LOGIC_VECTOR (27 downto 0) := "0000000000000110000000000001";
    constant ap_const_lv28_1FFE : STD_LOGIC_VECTOR (27 downto 0) := "0000000000000001111111111110";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';

    signal mul_res_V_fu_125_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal mul_res_V_reg_354 : STD_LOGIC_VECTOR (27 downto 0);
    signal ap_reg_ppstg_mul_res_V_reg_354_pp0_it1 : STD_LOGIC_VECTOR (27 downto 0);
    signal ap_reg_ppstg_mul_res_V_reg_354_pp0_it2 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_4_fu_147_p2 : STD_LOGIC_VECTOR (29 downto 0);
    signal r_V_4_reg_365 : STD_LOGIC_VECTOR (29 downto 0);
    signal r_V_10_fu_209_p2 : STD_LOGIC_VECTOR (36 downto 0);
    signal r_V_10_reg_370 : STD_LOGIC_VECTOR (36 downto 0);
    signal tmp_reg_375 : STD_LOGIC_VECTOR (13 downto 0);
    signal tmp_1_i_fu_327_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_1_i_reg_382 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_fu_83_p3 : STD_LOGIC_VECTOR (14 downto 0);
    signal r_V_1_fu_95_p3 : STD_LOGIC_VECTOR (25 downto 0);
    signal r_V_2_fu_107_p3 : STD_LOGIC_VECTOR (26 downto 0);
    signal r_V_2_cast_fu_115_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_cast_fu_91_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp1_fu_119_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_1_cast_fu_103_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal r_V_3_fu_131_p3 : STD_LOGIC_VECTOR (28 downto 0);
    signal rhs_V_cast_fu_143_p1 : STD_LOGIC_VECTOR (29 downto 0);
    signal lhs_V_cast_fu_139_p1 : STD_LOGIC_VECTOR (29 downto 0);
    signal r_V_5_fu_153_p3 : STD_LOGIC_VECTOR (31 downto 0);
    signal lhs_V_1_cast_fu_160_p1 : STD_LOGIC_VECTOR (32 downto 0);
    signal rhs_V_1_cast_fu_163_p1 : STD_LOGIC_VECTOR (32 downto 0);
    signal r_V_6_fu_167_p2 : STD_LOGIC_VECTOR (32 downto 0);
    signal r_V_7_fu_173_p3 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_V_2_cast_fu_180_p1 : STD_LOGIC_VECTOR (34 downto 0);
    signal rhs_V_2_cast_fu_184_p1 : STD_LOGIC_VECTOR (34 downto 0);
    signal r_V_8_fu_188_p2 : STD_LOGIC_VECTOR (34 downto 0);
    signal r_V_9_fu_194_p3 : STD_LOGIC_VECTOR (35 downto 0);
    signal lhs_V_3_cast_fu_201_p1 : STD_LOGIC_VECTOR (36 downto 0);
    signal rhs_V_3_cast_fu_205_p1 : STD_LOGIC_VECTOR (36 downto 0);
    signal r_V_11_fu_215_p3 : STD_LOGIC_VECTOR (37 downto 0);
    signal lhs_V_4_cast_fu_222_p1 : STD_LOGIC_VECTOR (38 downto 0);
    signal rhs_V_4_cast_fu_225_p1 : STD_LOGIC_VECTOR (38 downto 0);
    signal r_V_12_fu_229_p2 : STD_LOGIC_VECTOR (38 downto 0);
    signal r_V_13_fu_235_p3 : STD_LOGIC_VECTOR (39 downto 0);
    signal lhs_V_5_cast_fu_242_p1 : STD_LOGIC_VECTOR (40 downto 0);
    signal rhs_V_5_cast_fu_246_p1 : STD_LOGIC_VECTOR (40 downto 0);
    signal r_V_14_fu_250_p2 : STD_LOGIC_VECTOR (40 downto 0);
    signal r_V_15_fu_256_p3 : STD_LOGIC_VECTOR (41 downto 0);
    signal lhs_V_6_cast_fu_263_p1 : STD_LOGIC_VECTOR (42 downto 0);
    signal rhs_V_6_cast_fu_267_p1 : STD_LOGIC_VECTOR (42 downto 0);
    signal r_V_16_fu_271_p2 : STD_LOGIC_VECTOR (42 downto 0);
    signal phitmp_i_fu_287_p3 : STD_LOGIC_VECTOR (26 downto 0);
    signal phitmp2_i_fu_305_p3 : STD_LOGIC_VECTOR (14 downto 0);
    signal phitmp2_i_cast_fu_312_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal p_neg_i_fu_316_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal phitmp1_i_fu_298_p3 : STD_LOGIC_VECTOR (27 downto 0);
    signal p_neg1_i_fu_321_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal phitmp_i_cast_fu_294_p1 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_2_i_fu_333_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal p_i_fu_338_p2 : STD_LOGIC_VECTOR (27 downto 0);
    signal tmp_3_i_fu_343_p3 : STD_LOGIC_VECTOR (27 downto 0);


begin




    -- assign process. --
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_true = ap_true)) then
                ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(1) <= mul_res_V_reg_354(1);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(2) <= mul_res_V_reg_354(2);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(3) <= mul_res_V_reg_354(3);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(4) <= mul_res_V_reg_354(4);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(5) <= mul_res_V_reg_354(5);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(6) <= mul_res_V_reg_354(6);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(7) <= mul_res_V_reg_354(7);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(8) <= mul_res_V_reg_354(8);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(9) <= mul_res_V_reg_354(9);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(10) <= mul_res_V_reg_354(10);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(11) <= mul_res_V_reg_354(11);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(12) <= mul_res_V_reg_354(12);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(13) <= mul_res_V_reg_354(13);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(14) <= mul_res_V_reg_354(14);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(15) <= mul_res_V_reg_354(15);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(16) <= mul_res_V_reg_354(16);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(17) <= mul_res_V_reg_354(17);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(18) <= mul_res_V_reg_354(18);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(19) <= mul_res_V_reg_354(19);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(20) <= mul_res_V_reg_354(20);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(21) <= mul_res_V_reg_354(21);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(22) <= mul_res_V_reg_354(22);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(23) <= mul_res_V_reg_354(23);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(24) <= mul_res_V_reg_354(24);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(25) <= mul_res_V_reg_354(25);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(26) <= mul_res_V_reg_354(26);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(27) <= mul_res_V_reg_354(27);
                ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(1) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(1);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(2) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(2);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(3) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(3);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(4) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(4);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(5) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(5);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(6) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(6);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(7) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(7);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(8) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(8);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(9) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(9);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(10) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(10);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(11) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(11);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(12) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(12);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(13) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(13);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(14) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(14);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(15) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(15);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(16) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(16);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(17) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(17);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(18) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(18);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(19) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(19);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(20) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(20);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(21) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(21);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(22) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(22);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(23) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(23);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(24) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(24);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(25) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(25);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(26) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(26);
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(27) <= ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(27);
                mul_res_V_reg_354(1) <= mul_res_V_fu_125_p2(1);
    mul_res_V_reg_354(2) <= mul_res_V_fu_125_p2(2);
    mul_res_V_reg_354(3) <= mul_res_V_fu_125_p2(3);
    mul_res_V_reg_354(4) <= mul_res_V_fu_125_p2(4);
    mul_res_V_reg_354(5) <= mul_res_V_fu_125_p2(5);
    mul_res_V_reg_354(6) <= mul_res_V_fu_125_p2(6);
    mul_res_V_reg_354(7) <= mul_res_V_fu_125_p2(7);
    mul_res_V_reg_354(8) <= mul_res_V_fu_125_p2(8);
    mul_res_V_reg_354(9) <= mul_res_V_fu_125_p2(9);
    mul_res_V_reg_354(10) <= mul_res_V_fu_125_p2(10);
    mul_res_V_reg_354(11) <= mul_res_V_fu_125_p2(11);
    mul_res_V_reg_354(12) <= mul_res_V_fu_125_p2(12);
    mul_res_V_reg_354(13) <= mul_res_V_fu_125_p2(13);
    mul_res_V_reg_354(14) <= mul_res_V_fu_125_p2(14);
    mul_res_V_reg_354(15) <= mul_res_V_fu_125_p2(15);
    mul_res_V_reg_354(16) <= mul_res_V_fu_125_p2(16);
    mul_res_V_reg_354(17) <= mul_res_V_fu_125_p2(17);
    mul_res_V_reg_354(18) <= mul_res_V_fu_125_p2(18);
    mul_res_V_reg_354(19) <= mul_res_V_fu_125_p2(19);
    mul_res_V_reg_354(20) <= mul_res_V_fu_125_p2(20);
    mul_res_V_reg_354(21) <= mul_res_V_fu_125_p2(21);
    mul_res_V_reg_354(22) <= mul_res_V_fu_125_p2(22);
    mul_res_V_reg_354(23) <= mul_res_V_fu_125_p2(23);
    mul_res_V_reg_354(24) <= mul_res_V_fu_125_p2(24);
    mul_res_V_reg_354(25) <= mul_res_V_fu_125_p2(25);
    mul_res_V_reg_354(26) <= mul_res_V_fu_125_p2(26);
    mul_res_V_reg_354(27) <= mul_res_V_fu_125_p2(27);
                r_V_10_reg_370(1) <= r_V_10_fu_209_p2(1);
    r_V_10_reg_370(2) <= r_V_10_fu_209_p2(2);
    r_V_10_reg_370(3) <= r_V_10_fu_209_p2(3);
    r_V_10_reg_370(4) <= r_V_10_fu_209_p2(4);
    r_V_10_reg_370(5) <= r_V_10_fu_209_p2(5);
    r_V_10_reg_370(6) <= r_V_10_fu_209_p2(6);
    r_V_10_reg_370(7) <= r_V_10_fu_209_p2(7);
    r_V_10_reg_370(8) <= r_V_10_fu_209_p2(8);
    r_V_10_reg_370(9) <= r_V_10_fu_209_p2(9);
    r_V_10_reg_370(10) <= r_V_10_fu_209_p2(10);
    r_V_10_reg_370(11) <= r_V_10_fu_209_p2(11);
    r_V_10_reg_370(12) <= r_V_10_fu_209_p2(12);
    r_V_10_reg_370(13) <= r_V_10_fu_209_p2(13);
    r_V_10_reg_370(14) <= r_V_10_fu_209_p2(14);
    r_V_10_reg_370(15) <= r_V_10_fu_209_p2(15);
    r_V_10_reg_370(16) <= r_V_10_fu_209_p2(16);
    r_V_10_reg_370(17) <= r_V_10_fu_209_p2(17);
    r_V_10_reg_370(18) <= r_V_10_fu_209_p2(18);
    r_V_10_reg_370(19) <= r_V_10_fu_209_p2(19);
    r_V_10_reg_370(20) <= r_V_10_fu_209_p2(20);
    r_V_10_reg_370(21) <= r_V_10_fu_209_p2(21);
    r_V_10_reg_370(22) <= r_V_10_fu_209_p2(22);
    r_V_10_reg_370(23) <= r_V_10_fu_209_p2(23);
    r_V_10_reg_370(24) <= r_V_10_fu_209_p2(24);
    r_V_10_reg_370(25) <= r_V_10_fu_209_p2(25);
    r_V_10_reg_370(26) <= r_V_10_fu_209_p2(26);
    r_V_10_reg_370(27) <= r_V_10_fu_209_p2(27);
    r_V_10_reg_370(28) <= r_V_10_fu_209_p2(28);
    r_V_10_reg_370(29) <= r_V_10_fu_209_p2(29);
    r_V_10_reg_370(30) <= r_V_10_fu_209_p2(30);
    r_V_10_reg_370(31) <= r_V_10_fu_209_p2(31);
    r_V_10_reg_370(32) <= r_V_10_fu_209_p2(32);
    r_V_10_reg_370(33) <= r_V_10_fu_209_p2(33);
    r_V_10_reg_370(34) <= r_V_10_fu_209_p2(34);
    r_V_10_reg_370(35) <= r_V_10_fu_209_p2(35);
    r_V_10_reg_370(36) <= r_V_10_fu_209_p2(36);
                r_V_4_reg_365(1) <= r_V_4_fu_147_p2(1);
    r_V_4_reg_365(2) <= r_V_4_fu_147_p2(2);
    r_V_4_reg_365(3) <= r_V_4_fu_147_p2(3);
    r_V_4_reg_365(4) <= r_V_4_fu_147_p2(4);
    r_V_4_reg_365(5) <= r_V_4_fu_147_p2(5);
    r_V_4_reg_365(6) <= r_V_4_fu_147_p2(6);
    r_V_4_reg_365(7) <= r_V_4_fu_147_p2(7);
    r_V_4_reg_365(8) <= r_V_4_fu_147_p2(8);
    r_V_4_reg_365(9) <= r_V_4_fu_147_p2(9);
    r_V_4_reg_365(10) <= r_V_4_fu_147_p2(10);
    r_V_4_reg_365(11) <= r_V_4_fu_147_p2(11);
    r_V_4_reg_365(12) <= r_V_4_fu_147_p2(12);
    r_V_4_reg_365(13) <= r_V_4_fu_147_p2(13);
    r_V_4_reg_365(14) <= r_V_4_fu_147_p2(14);
    r_V_4_reg_365(15) <= r_V_4_fu_147_p2(15);
    r_V_4_reg_365(16) <= r_V_4_fu_147_p2(16);
    r_V_4_reg_365(17) <= r_V_4_fu_147_p2(17);
    r_V_4_reg_365(18) <= r_V_4_fu_147_p2(18);
    r_V_4_reg_365(19) <= r_V_4_fu_147_p2(19);
    r_V_4_reg_365(20) <= r_V_4_fu_147_p2(20);
    r_V_4_reg_365(21) <= r_V_4_fu_147_p2(21);
    r_V_4_reg_365(22) <= r_V_4_fu_147_p2(22);
    r_V_4_reg_365(23) <= r_V_4_fu_147_p2(23);
    r_V_4_reg_365(24) <= r_V_4_fu_147_p2(24);
    r_V_4_reg_365(25) <= r_V_4_fu_147_p2(25);
    r_V_4_reg_365(26) <= r_V_4_fu_147_p2(26);
    r_V_4_reg_365(27) <= r_V_4_fu_147_p2(27);
    r_V_4_reg_365(28) <= r_V_4_fu_147_p2(28);
    r_V_4_reg_365(29) <= r_V_4_fu_147_p2(29);
                tmp_1_i_reg_382(1) <= tmp_1_i_fu_327_p2(1);
    tmp_1_i_reg_382(2) <= tmp_1_i_fu_327_p2(2);
    tmp_1_i_reg_382(3) <= tmp_1_i_fu_327_p2(3);
    tmp_1_i_reg_382(4) <= tmp_1_i_fu_327_p2(4);
    tmp_1_i_reg_382(5) <= tmp_1_i_fu_327_p2(5);
    tmp_1_i_reg_382(6) <= tmp_1_i_fu_327_p2(6);
    tmp_1_i_reg_382(7) <= tmp_1_i_fu_327_p2(7);
    tmp_1_i_reg_382(8) <= tmp_1_i_fu_327_p2(8);
    tmp_1_i_reg_382(9) <= tmp_1_i_fu_327_p2(9);
    tmp_1_i_reg_382(10) <= tmp_1_i_fu_327_p2(10);
    tmp_1_i_reg_382(11) <= tmp_1_i_fu_327_p2(11);
    tmp_1_i_reg_382(12) <= tmp_1_i_fu_327_p2(12);
    tmp_1_i_reg_382(13) <= tmp_1_i_fu_327_p2(13);
    tmp_1_i_reg_382(14) <= tmp_1_i_fu_327_p2(14);
    tmp_1_i_reg_382(15) <= tmp_1_i_fu_327_p2(15);
    tmp_1_i_reg_382(16) <= tmp_1_i_fu_327_p2(16);
    tmp_1_i_reg_382(17) <= tmp_1_i_fu_327_p2(17);
    tmp_1_i_reg_382(18) <= tmp_1_i_fu_327_p2(18);
    tmp_1_i_reg_382(19) <= tmp_1_i_fu_327_p2(19);
    tmp_1_i_reg_382(20) <= tmp_1_i_fu_327_p2(20);
    tmp_1_i_reg_382(21) <= tmp_1_i_fu_327_p2(21);
    tmp_1_i_reg_382(22) <= tmp_1_i_fu_327_p2(22);
    tmp_1_i_reg_382(23) <= tmp_1_i_fu_327_p2(23);
    tmp_1_i_reg_382(24) <= tmp_1_i_fu_327_p2(24);
    tmp_1_i_reg_382(25) <= tmp_1_i_fu_327_p2(25);
    tmp_1_i_reg_382(26) <= tmp_1_i_fu_327_p2(26);
    tmp_1_i_reg_382(27) <= tmp_1_i_fu_327_p2(27);
                tmp_reg_375 <= r_V_16_fu_271_p2(42 downto 29);
            end if;
        end if;
    end process;
    mul_res_V_reg_354(0) <= '0';
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it1(0) <= '0';
    ap_reg_ppstg_mul_res_V_reg_354_pp0_it2(0) <= '0';
    r_V_4_reg_365(0) <= '0';
    r_V_10_reg_370(0) <= '0';
    tmp_1_i_reg_382(0) <= '0';
    ap_return <= tmp_3_i_fu_343_p3(15 - 1 downto 0);
    lhs_V_1_cast_fu_160_p1 <= std_logic_vector(resize(unsigned(r_V_4_reg_365),33));
    lhs_V_2_cast_fu_180_p1 <= std_logic_vector(resize(unsigned(r_V_6_fu_167_p2),35));
    lhs_V_3_cast_fu_201_p1 <= std_logic_vector(resize(unsigned(r_V_8_fu_188_p2),37));
    lhs_V_4_cast_fu_222_p1 <= std_logic_vector(resize(unsigned(r_V_10_reg_370),39));
    lhs_V_5_cast_fu_242_p1 <= std_logic_vector(resize(unsigned(r_V_12_fu_229_p2),41));
    lhs_V_6_cast_fu_263_p1 <= std_logic_vector(resize(unsigned(r_V_14_fu_250_p2),43));
    lhs_V_cast_fu_139_p1 <= std_logic_vector(resize(unsigned(mul_res_V_fu_125_p2),30));
    mul_res_V_fu_125_p2 <= std_logic_vector(unsigned(tmp1_fu_119_p2) + unsigned(r_V_1_cast_fu_103_p1));
    p_i_fu_338_p2 <= std_logic_vector(unsigned(tmp_1_i_reg_382) + unsigned(ap_const_lv28_1FFE));
    p_neg1_i_fu_321_p2 <= std_logic_vector(unsigned(p_neg_i_fu_316_p2) - unsigned(phitmp1_i_fu_298_p3));
    p_neg_i_fu_316_p2 <= std_logic_vector(unsigned(ap_reg_ppstg_mul_res_V_reg_354_pp0_it2) - unsigned(phitmp2_i_cast_fu_312_p1));
    phitmp1_i_fu_298_p3 <= (tmp_reg_375 & ap_const_lv14_0);
    phitmp2_i_cast_fu_312_p1 <= std_logic_vector(resize(unsigned(phitmp2_i_fu_305_p3),28));
    phitmp2_i_fu_305_p3 <= (tmp_reg_375 & ap_const_lv1_0);
    phitmp_i_cast_fu_294_p1 <= std_logic_vector(resize(unsigned(phitmp_i_fu_287_p3),28));
    phitmp_i_fu_287_p3 <= (tmp_reg_375 & ap_const_lv13_0);
    r_V_10_fu_209_p2 <= std_logic_vector(unsigned(lhs_V_3_cast_fu_201_p1) + unsigned(rhs_V_3_cast_fu_205_p1));
    r_V_11_fu_215_p3 <= (ap_reg_ppstg_mul_res_V_reg_354_pp0_it1 & ap_const_lv10_0);
    r_V_12_fu_229_p2 <= std_logic_vector(unsigned(lhs_V_4_cast_fu_222_p1) + unsigned(rhs_V_4_cast_fu_225_p1));
    r_V_13_fu_235_p3 <= (ap_reg_ppstg_mul_res_V_reg_354_pp0_it1 & ap_const_lv12_0);
    r_V_14_fu_250_p2 <= std_logic_vector(unsigned(lhs_V_5_cast_fu_242_p1) + unsigned(rhs_V_5_cast_fu_246_p1));
    r_V_15_fu_256_p3 <= (ap_reg_ppstg_mul_res_V_reg_354_pp0_it1 & ap_const_lv14_0);
    r_V_16_fu_271_p2 <= std_logic_vector(unsigned(lhs_V_6_cast_fu_263_p1) + unsigned(rhs_V_6_cast_fu_267_p1));
    r_V_1_cast_fu_103_p1 <= std_logic_vector(resize(unsigned(r_V_1_fu_95_p3),28));
    r_V_1_fu_95_p3 <= (data_in_V & ap_const_lv12_0);
    r_V_2_cast_fu_115_p1 <= std_logic_vector(resize(unsigned(r_V_2_fu_107_p3),28));
    r_V_2_fu_107_p3 <= (data_in_V & ap_const_lv13_0);
    r_V_3_fu_131_p3 <= (mul_res_V_fu_125_p2 & ap_const_lv1_0);
    r_V_4_fu_147_p2 <= std_logic_vector(unsigned(rhs_V_cast_fu_143_p1) + unsigned(lhs_V_cast_fu_139_p1));
    r_V_5_fu_153_p3 <= (mul_res_V_reg_354 & ap_const_lv4_0);
    r_V_6_fu_167_p2 <= std_logic_vector(unsigned(lhs_V_1_cast_fu_160_p1) + unsigned(rhs_V_1_cast_fu_163_p1));
    r_V_7_fu_173_p3 <= (mul_res_V_reg_354 & ap_const_lv6_0);
    r_V_8_fu_188_p2 <= std_logic_vector(unsigned(lhs_V_2_cast_fu_180_p1) + unsigned(rhs_V_2_cast_fu_184_p1));
    r_V_9_fu_194_p3 <= (mul_res_V_reg_354 & ap_const_lv8_0);
    r_V_cast_fu_91_p1 <= std_logic_vector(resize(unsigned(r_V_fu_83_p3),28));
    r_V_fu_83_p3 <= (data_in_V & ap_const_lv1_0);
    rhs_V_1_cast_fu_163_p1 <= std_logic_vector(resize(unsigned(r_V_5_fu_153_p3),33));
    rhs_V_2_cast_fu_184_p1 <= std_logic_vector(resize(unsigned(r_V_7_fu_173_p3),35));
    rhs_V_3_cast_fu_205_p1 <= std_logic_vector(resize(unsigned(r_V_9_fu_194_p3),37));
    rhs_V_4_cast_fu_225_p1 <= std_logic_vector(resize(unsigned(r_V_11_fu_215_p3),39));
    rhs_V_5_cast_fu_246_p1 <= std_logic_vector(resize(unsigned(r_V_13_fu_235_p3),41));
    rhs_V_6_cast_fu_267_p1 <= std_logic_vector(resize(unsigned(r_V_15_fu_256_p3),43));
    rhs_V_cast_fu_143_p1 <= std_logic_vector(resize(unsigned(r_V_3_fu_131_p3),30));
    tmp1_fu_119_p2 <= std_logic_vector(unsigned(r_V_2_cast_fu_115_p1) + unsigned(r_V_cast_fu_91_p1));
    tmp_1_i_fu_327_p2 <= std_logic_vector(unsigned(p_neg1_i_fu_321_p2) - unsigned(phitmp_i_cast_fu_294_p1));
    tmp_2_i_fu_333_p2 <= "1" when (unsigned(tmp_1_i_reg_382) > unsigned(ap_const_lv28_6001)) else "0";
    tmp_3_i_fu_343_p3 <= 
        p_i_fu_338_p2 when (tmp_2_i_fu_333_p2(0) = '1') else 
        tmp_1_i_reg_382;
end behav;
