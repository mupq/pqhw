--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/

-- TestBench Template 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


entity rejection_module_tb is
  generic (
    RAM_DEPTH        : integer               := 64;
    NUMBER_OF_BLOCKS : integer               := 16;
    --------------------------General -----------------------------------------
    N_ELEMENTS       : integer               := 512;
    PRIME_P_WIDTH    : integer               := 14;
    PRIME_P          : unsigned              := to_unsigned(12289, 14);
    -----------------------  Sparse Mul Core ----------------------------------
    KAPPA            : integer               := 23;
    HASH_BLOCKS      : integer               := 4;
    HASH_WIDTH       : integer               := 64;
    --------------------------General --------------------------------------
    ZETA             : unsigned              := to_unsigned(6145, 13);
    D_BLISS          : integer               := 10;
    MODULUS_P_BLISS  : unsigned              := to_unsigned(24, 5);
    -----------------------  Sparse Mul Core ------------------------------------------
    CORES            : integer               := 8;
    WIDTH_S1         : integer               := 2;
    WIDTH_S2         : integer               := 3;
    --Used to initialize the right s (s1 or s2)
    INIT_TABLE       : integer               := 0;
    c_delay          : integer range 0 to 16 := 2;
    ---------------------------------------------------------------------------
    MAX_RES_WIDTH    : integer               := 6
    );
  port (
    error_happened_out    : out std_logic := '0';
    end_of_simulation_out : out std_logic := '0'
    );
end rejection_module_tb;

architecture behavior of rejection_module_tb is
  signal end_of_simulation : std_logic := '0';
  signal error_happened    : std_logic := '0';


  signal   clk           : std_logic;
  constant clk_period    : time    := 10 ns;
  signal   cycle_counter : integer := 0;
  type     ram_type is array (0 to N_ELEMENTS-1) of signed(32-1 downto 0);


  signal y1 : ram_type := (to_signed(110,32), to_signed(12250,32), to_signed(12096,32), to_signed(209,32), to_signed(7,32), to_signed(12282,32), to_signed(12131,32), to_signed(97,32), to_signed(142,32), to_signed(12210,32), to_signed(115,32), to_signed(12113,32), to_signed(12005,32), to_signed(253,32), to_signed(209,32), to_signed(231,32), to_signed(12047,32), to_signed(12259,32), to_signed(12145,32), to_signed(254,32), to_signed(47,32), to_signed(15,32), to_signed(12271,32), to_signed(251,32), to_signed(282,32), to_signed(12173,32), to_signed(12121,32), to_signed(28,32), to_signed(12061,32), to_signed(11930,32), to_signed(12191,32), to_signed(177,32), to_signed(214,32), to_signed(12162,32), to_signed(12225,32), to_signed(50,32), to_signed(12237,32), to_signed(11921,32), to_signed(168,32), to_signed(11910,32), to_signed(310,32), to_signed(11785,32), to_signed(12281,32), to_signed(12061,32), to_signed(69,32), to_signed(12182,32), to_signed(12285,32), to_signed(12020,32), to_signed(267,32), to_signed(12029,32), to_signed(220,32), to_signed(364,32), to_signed(12233,32), to_signed(12202,32), to_signed(171,32), to_signed(12140,32), to_signed(208,32), to_signed(23,32), to_signed(668,32), to_signed(11948,32), to_signed(70,32), to_signed(70,32), to_signed(187,32), to_signed(12219,32), to_signed(12090,32), to_signed(12195,32), to_signed(38,32), to_signed(12084,32), to_signed(12271,32), to_signed(85,32), to_signed(117,32), to_signed(12237,32), to_signed(12264,32), to_signed(11887,32), to_signed(295,32), to_signed(12121,32), to_signed(71,32), to_signed(11977,32), to_signed(12013,32), to_signed(65,32), to_signed(212,32), to_signed(282,32), to_signed(340,32), to_signed(0,32), to_signed(12150,32), to_signed(11953,32), to_signed(12180,32), to_signed(28,32), to_signed(12054,32), to_signed(34,32), to_signed(12208,32), to_signed(56,32), to_signed(11985,32), to_signed(12240,32), to_signed(12213,32), to_signed(111,32), to_signed(11782,32), to_signed(96,32), to_signed(12226,32), to_signed(230,32), to_signed(310,32), to_signed(19,32), to_signed(172,32), to_signed(12037,32), to_signed(69,32), to_signed(12021,32), to_signed(12246,32), to_signed(12234,32), to_signed(11985,32), to_signed(23,32), to_signed(12175,32), to_signed(12234,32), to_signed(282,32), to_signed(232,32), to_signed(12216,32), to_signed(61,32), to_signed(12183,32), to_signed(12136,32), to_signed(147,32), to_signed(12279,32), to_signed(11928,32), to_signed(12195,32), to_signed(245,32), to_signed(108,32), to_signed(155,32), to_signed(11801,32), to_signed(11945,32), to_signed(12154,32), to_signed(12141,32), to_signed(11889,32), to_signed(94,32), to_signed(78,32), to_signed(11979,32), to_signed(4,32), to_signed(12244,32), to_signed(12159,32), to_signed(12131,32), to_signed(12082,32), to_signed(12151,32), to_signed(101,32), to_signed(8,32), to_signed(12058,32), to_signed(45,32), to_signed(23,32), to_signed(143,32), to_signed(50,32), to_signed(125,32), to_signed(292,32), to_signed(12219,32), to_signed(196,32), to_signed(12116,32), to_signed(60,32), to_signed(248,32), to_signed(111,32), to_signed(171,32), to_signed(12162,32), to_signed(12239,32), to_signed(12190,32), to_signed(12081,32), to_signed(12058,32), to_signed(12242,32), to_signed(11956,32), to_signed(11980,32), to_signed(143,32), to_signed(12263,32), to_signed(12196,32), to_signed(12155,32), to_signed(112,32), to_signed(11944,32), to_signed(80,32), to_signed(492,32), to_signed(11970,32), to_signed(41,32), to_signed(271,32), to_signed(49,32), to_signed(96,32), to_signed(12029,32), to_signed(12010,32), to_signed(226,32), to_signed(239,32), to_signed(353,32), to_signed(104,32), to_signed(59,32), to_signed(12063,32), to_signed(274,32), to_signed(82,32), to_signed(12259,32), to_signed(260,32), to_signed(394,32), to_signed(11692,32), to_signed(414,32), to_signed(11904,32), to_signed(12137,32), to_signed(129,32), to_signed(11765,32), to_signed(12041,32), to_signed(1,32), to_signed(12150,32), to_signed(3,32), to_signed(501,32), to_signed(12192,32), to_signed(12172,32), to_signed(287,32), to_signed(12137,32), to_signed(12249,32), to_signed(12182,32), to_signed(12239,32), to_signed(29,32), to_signed(12176,32), to_signed(12257,32), to_signed(12005,32), to_signed(12256,32), to_signed(190,32), to_signed(12231,32), to_signed(12259,32), to_signed(12122,32), to_signed(288,32), to_signed(5,32), to_signed(168,32), to_signed(111,32), to_signed(86,32), to_signed(12074,32), to_signed(12282,32), to_signed(11905,32), to_signed(9,32), to_signed(12166,32), to_signed(181,32), to_signed(11871,32), to_signed(57,32), to_signed(44,32), to_signed(12110,32), to_signed(12114,32), to_signed(34,32), to_signed(398,32), to_signed(24,32), to_signed(111,32), to_signed(258,32), to_signed(11996,32), to_signed(1,32), to_signed(226,32), to_signed(234,32), to_signed(302,32), to_signed(12235,32), to_signed(377,32), to_signed(12197,32), to_signed(12261,32), to_signed(12169,32), to_signed(6,32), to_signed(475,32), to_signed(59,32), to_signed(137,32), to_signed(12108,32), to_signed(10,32), to_signed(12138,32), to_signed(41,32), to_signed(199,32), to_signed(12160,32), to_signed(329,32), to_signed(12233,32), to_signed(163,32), to_signed(12232,32), to_signed(211,32), to_signed(12275,32), to_signed(12230,32), to_signed(12075,32), to_signed(68,32), to_signed(12171,32), to_signed(12044,32), to_signed(280,32), to_signed(192,32), to_signed(12222,32), to_signed(12169,32), to_signed(439,32), to_signed(277,32), to_signed(12235,32), to_signed(12045,32), to_signed(311,32), to_signed(12175,32), to_signed(433,32), to_signed(12137,32), to_signed(16,32), to_signed(36,32), to_signed(163,32), to_signed(12277,32), to_signed(11827,32), to_signed(12287,32), to_signed(12267,32), to_signed(12284,32), to_signed(12213,32), to_signed(11866,32), to_signed(144,32), to_signed(12228,32), to_signed(12165,32), to_signed(15,32), to_signed(188,32), to_signed(0,32), to_signed(12263,32), to_signed(11901,32), to_signed(36,32), to_signed(39,32), to_signed(12009,32), to_signed(12160,32), to_signed(12086,32), to_signed(12123,32), to_signed(432,32), to_signed(12078,32), to_signed(12171,32), to_signed(365,32), to_signed(130,32), to_signed(12241,32), to_signed(180,32), to_signed(121,32), to_signed(390,32), to_signed(12144,32), to_signed(134,32), to_signed(12257,32), to_signed(12237,32), to_signed(204,32), to_signed(122,32), to_signed(12279,32), to_signed(11754,32), to_signed(190,32), to_signed(225,32), to_signed(11977,32), to_signed(12167,32), to_signed(47,32), to_signed(12183,32), to_signed(363,32), to_signed(17,32), to_signed(12258,32), to_signed(11966,32), to_signed(12265,32), to_signed(93,32), to_signed(11982,32), to_signed(241,32), to_signed(12043,32), to_signed(12007,32), to_signed(415,32), to_signed(12217,32), to_signed(12276,32), to_signed(304,32), to_signed(12281,32), to_signed(12050,32), to_signed(104,32), to_signed(11968,32), to_signed(193,32), to_signed(86,32), to_signed(220,32), to_signed(242,32), to_signed(12009,32), to_signed(12249,32), to_signed(69,32), to_signed(303,32), to_signed(12064,32), to_signed(46,32), to_signed(78,32), to_signed(169,32), to_signed(182,32), to_signed(12221,32), to_signed(11899,32), to_signed(251,32), to_signed(12280,32), to_signed(12161,32), to_signed(11912,32), to_signed(12047,32), to_signed(424,32), to_signed(12164,32), to_signed(12047,32), to_signed(150,32), to_signed(12176,32), to_signed(12225,32), to_signed(12181,32), to_signed(181,32), to_signed(12092,32), to_signed(12252,32), to_signed(12115,32), to_signed(12163,32), to_signed(135,32), to_signed(422,32), to_signed(126,32), to_signed(11726,32), to_signed(151,32), to_signed(27,32), to_signed(12082,32), to_signed(12018,32), to_signed(269,32), to_signed(408,32), to_signed(110,32), to_signed(305,32), to_signed(513,32), to_signed(12161,32), to_signed(12155,32), to_signed(305,32), to_signed(171,32), to_signed(64,32), to_signed(47,32), to_signed(12195,32), to_signed(202,32), to_signed(12041,32), to_signed(12184,32), to_signed(12067,32), to_signed(97,32), to_signed(12050,32), to_signed(11999,32), to_signed(161,32), to_signed(11775,32), to_signed(330,32), to_signed(492,32), to_signed(12053,32), to_signed(280,32), to_signed(175,32), to_signed(32,32), to_signed(12051,32), to_signed(39,32), to_signed(12133,32), to_signed(23,32), to_signed(208,32), to_signed(12266,32), to_signed(12121,32), to_signed(11942,32), to_signed(226,32), to_signed(12039,32), to_signed(11806,32), to_signed(292,32), to_signed(12056,32), to_signed(12147,32), to_signed(149,32), to_signed(33,32), to_signed(12087,32), to_signed(12237,32), to_signed(12061,32), to_signed(293,32), to_signed(12247,32), to_signed(11904,32), to_signed(11913,32), to_signed(54,32), to_signed(11787,32), to_signed(12256,32), to_signed(324,32), to_signed(18,32), to_signed(11827,32), to_signed(206,32), to_signed(26,32), to_signed(12001,32), to_signed(192,32), to_signed(249,32), to_signed(116,32), to_signed(232,32), to_signed(136,32), to_signed(294,32), to_signed(12185,32), to_signed(19,32), to_signed(340,32), to_signed(12111,32), to_signed(358,32), to_signed(85,32), to_signed(126,32), to_signed(35,32), to_signed(12113,32), to_signed(197,32), to_signed(12185,32), to_signed(12272,32), to_signed(623,32), to_signed(301,32), to_signed(12235,32), to_signed(2,32), to_signed(11872,32), to_signed(126,32), to_signed(11767,32), to_signed(12226,32), to_signed(12099,32), to_signed(311,32), to_signed(6,32), to_signed(12269,32), to_signed(12154,32), to_signed(12146,32), to_signed(11975,32), to_signed(12258,32), to_signed(125,32), to_signed(92,32), to_signed(11819,32), to_signed(12256,32), to_signed(341,32), to_signed(161,32), to_signed(12209,32), to_signed(57,32), to_signed(242,32), to_signed(268,32), to_signed(12251,32), to_signed(26,32), to_signed(11950,32), to_signed(12260,32), to_signed(12219,32), to_signed(12122,32), to_signed(253,32), to_signed(12208,32), to_signed(124,32), to_signed(12187,32), to_signed(155,32), to_signed(12128,32), to_signed(52,32), to_signed(12248,32), to_signed(11757,32), to_signed(438,32), to_signed(320,32), to_signed(12165,32), to_signed(277,32), to_signed(12071,32), to_signed(12062,32), to_signed(12267,32), to_signed(163,32), to_signed(37,32));


  signal y2 : ram_type := (to_signed(284,32), to_signed(12174,32), to_signed(0,32), to_signed(55,32), to_signed(12096,32), to_signed(12207,32), to_signed(299,32), to_signed(12152,32), to_signed(12027,32), to_signed(12227,32), to_signed(12223,32), to_signed(12031,32), to_signed(12189,32), to_signed(12264,32), to_signed(12274,32), to_signed(12001,32), to_signed(11960,32), to_signed(12170,32), to_signed(12205,32), to_signed(637,32), to_signed(12285,32), to_signed(12123,32), to_signed(12025,32), to_signed(12015,32), to_signed(121,32), to_signed(12173,32), to_signed(12182,32), to_signed(65,32), to_signed(12243,32), to_signed(12173,32), to_signed(11956,32), to_signed(198,32), to_signed(11856,32), to_signed(83,32), to_signed(12271,32), to_signed(11902,32), to_signed(376,32), to_signed(350,32), to_signed(77,32), to_signed(128,32), to_signed(12041,32), to_signed(182,32), to_signed(242,32), to_signed(12287,32), to_signed(149,32), to_signed(12227,32), to_signed(12273,32), to_signed(12281,32), to_signed(11885,32), to_signed(12042,32), to_signed(12189,32), to_signed(210,32), to_signed(410,32), to_signed(193,32), to_signed(231,32), to_signed(12286,32), to_signed(11985,32), to_signed(174,32), to_signed(12175,32), to_signed(12022,32), to_signed(12242,32), to_signed(12186,32), to_signed(276,32), to_signed(12135,32), to_signed(236,32), to_signed(25,32), to_signed(12034,32), to_signed(324,32), to_signed(342,32), to_signed(12279,32), to_signed(12174,32), to_signed(11839,32), to_signed(11978,32), to_signed(12143,32), to_signed(43,32), to_signed(97,32), to_signed(37,32), to_signed(12287,32), to_signed(74,32), to_signed(12249,32), to_signed(12203,32), to_signed(346,32), to_signed(12226,32), to_signed(222,32), to_signed(12170,32), to_signed(12004,32), to_signed(402,32), to_signed(12251,32), to_signed(11795,32), to_signed(327,32), to_signed(166,32), to_signed(12265,32), to_signed(12157,32), to_signed(12082,32), to_signed(1,32), to_signed(12,32), to_signed(403,32), to_signed(12153,32), to_signed(23,32), to_signed(12208,32), to_signed(584,32), to_signed(328,32), to_signed(12079,32), to_signed(12121,32), to_signed(80,32), to_signed(12049,32), to_signed(12202,32), to_signed(12168,32), to_signed(12158,32), to_signed(12260,32), to_signed(64,32), to_signed(81,32), to_signed(12245,32), to_signed(12246,32), to_signed(12284,32), to_signed(12286,32), to_signed(11962,32), to_signed(94,32), to_signed(12261,32), to_signed(12074,32), to_signed(12033,32), to_signed(8,32), to_signed(12134,32), to_signed(26,32), to_signed(12144,32), to_signed(117,32), to_signed(12158,32), to_signed(12231,32), to_signed(20,32), to_signed(129,32), to_signed(12116,32), to_signed(12142,32), to_signed(12112,32), to_signed(12248,32), to_signed(76,32), to_signed(11962,32), to_signed(281,32), to_signed(12123,32), to_signed(168,32), to_signed(12200,32), to_signed(2,32), to_signed(406,32), to_signed(363,32), to_signed(12151,32), to_signed(256,32), to_signed(12187,32), to_signed(110,32), to_signed(11980,32), to_signed(11933,32), to_signed(12082,32), to_signed(49,32), to_signed(12019,32), to_signed(11799,32), to_signed(71,32), to_signed(12210,32), to_signed(334,32), to_signed(12271,32), to_signed(12011,32), to_signed(201,32), to_signed(12096,32), to_signed(80,32), to_signed(68,32), to_signed(133,32), to_signed(108,32), to_signed(59,32), to_signed(213,32), to_signed(12061,32), to_signed(91,32), to_signed(12089,32), to_signed(12203,32), to_signed(12209,32), to_signed(117,32), to_signed(233,32), to_signed(11986,32), to_signed(12224,32), to_signed(12158,32), to_signed(72,32), to_signed(38,32), to_signed(12178,32), to_signed(405,32), to_signed(158,32), to_signed(12262,32), to_signed(12126,32), to_signed(12183,32), to_signed(12125,32), to_signed(470,32), to_signed(151,32), to_signed(175,32), to_signed(12224,32), to_signed(85,32), to_signed(103,32), to_signed(12239,32), to_signed(123,32), to_signed(239,32), to_signed(104,32), to_signed(12157,32), to_signed(12257,32), to_signed(12221,32), to_signed(56,32), to_signed(12227,32), to_signed(12203,32), to_signed(110,32), to_signed(11954,32), to_signed(11860,32), to_signed(12044,32), to_signed(12208,32), to_signed(10,32), to_signed(12209,32), to_signed(173,32), to_signed(107,32), to_signed(320,32), to_signed(18,32), to_signed(40,32), to_signed(244,32), to_signed(12198,32), to_signed(12065,32), to_signed(12250,32), to_signed(2,32), to_signed(83,32), to_signed(12178,32), to_signed(12097,32), to_signed(12153,32), to_signed(166,32), to_signed(12144,32), to_signed(242,32), to_signed(12076,32), to_signed(11894,32), to_signed(12283,32), to_signed(11829,32), to_signed(59,32), to_signed(12181,32), to_signed(11966,32), to_signed(12150,32), to_signed(23,32), to_signed(11986,32), to_signed(130,32), to_signed(12250,32), to_signed(42,32), to_signed(98,32), to_signed(72,32), to_signed(136,32), to_signed(12180,32), to_signed(86,32), to_signed(12183,32), to_signed(193,32), to_signed(11917,32), to_signed(12179,32), to_signed(11806,32), to_signed(12209,32), to_signed(12062,32), to_signed(266,32), to_signed(12085,32), to_signed(14,32), to_signed(12204,32), to_signed(53,32), to_signed(12201,32), to_signed(12077,32), to_signed(12234,32), to_signed(89,32), to_signed(425,32), to_signed(111,32), to_signed(119,32), to_signed(12086,32), to_signed(134,32), to_signed(354,32), to_signed(12088,32), to_signed(128,32), to_signed(367,32), to_signed(12168,32), to_signed(76,32), to_signed(203,32), to_signed(12056,32), to_signed(12022,32), to_signed(12005,32), to_signed(169,32), to_signed(12127,32), to_signed(11991,32), to_signed(182,32), to_signed(73,32), to_signed(12190,32), to_signed(182,32), to_signed(87,32), to_signed(12166,32), to_signed(194,32), to_signed(628,32), to_signed(12236,32), to_signed(12214,32), to_signed(110,32), to_signed(12115,32), to_signed(12207,32), to_signed(11949,32), to_signed(12101,32), to_signed(12153,32), to_signed(12066,32), to_signed(12170,32), to_signed(12079,32), to_signed(12284,32), to_signed(12,32), to_signed(141,32), to_signed(11905,32), to_signed(12160,32), to_signed(141,32), to_signed(12249,32), to_signed(12009,32), to_signed(12048,32), to_signed(11977,32), to_signed(12180,32), to_signed(272,32), to_signed(472,32), to_signed(116,32), to_signed(12260,32), to_signed(174,32), to_signed(195,32), to_signed(48,32), to_signed(285,32), to_signed(281,32), to_signed(372,32), to_signed(12216,32), to_signed(11930,32), to_signed(148,32), to_signed(450,32), to_signed(283,32), to_signed(12085,32), to_signed(12167,32), to_signed(12053,32), to_signed(12053,32), to_signed(11934,32), to_signed(430,32), to_signed(11879,32), to_signed(123,32), to_signed(12284,32), to_signed(103,32), to_signed(7,32), to_signed(74,32), to_signed(229,32), to_signed(12070,32), to_signed(12204,32), to_signed(12105,32), to_signed(263,32), to_signed(235,32), to_signed(178,32), to_signed(12018,32), to_signed(156,32), to_signed(104,32), to_signed(12057,32), to_signed(139,32), to_signed(12208,32), to_signed(12174,32), to_signed(183,32), to_signed(12103,32), to_signed(12141,32), to_signed(12284,32), to_signed(11916,32), to_signed(11978,32), to_signed(12140,32), to_signed(81,32), to_signed(193,32), to_signed(12170,32), to_signed(12141,32), to_signed(12132,32), to_signed(12190,32), to_signed(12061,32), to_signed(42,32), to_signed(111,32), to_signed(12253,32), to_signed(229,32), to_signed(165,32), to_signed(12035,32), to_signed(57,32), to_signed(278,32), to_signed(90,32), to_signed(12086,32), to_signed(279,32), to_signed(324,32), to_signed(245,32), to_signed(169,32), to_signed(12241,32), to_signed(240,32), to_signed(327,32), to_signed(385,32), to_signed(12112,32), to_signed(80,32), to_signed(34,32), to_signed(429,32), to_signed(12272,32), to_signed(293,32), to_signed(12058,32), to_signed(176,32), to_signed(12274,32), to_signed(12109,32), to_signed(12183,32), to_signed(9,32), to_signed(283,32), to_signed(12020,32), to_signed(221,32), to_signed(93,32), to_signed(471,32), to_signed(178,32), to_signed(12243,32), to_signed(56,32), to_signed(12145,32), to_signed(149,32), to_signed(20,32), to_signed(22,32), to_signed(202,32), to_signed(12206,32), to_signed(120,32), to_signed(258,32), to_signed(27,32), to_signed(12209,32), to_signed(12148,32), to_signed(11894,32), to_signed(12160,32), to_signed(104,32), to_signed(138,32), to_signed(23,32), to_signed(12255,32), to_signed(12103,32), to_signed(12229,32), to_signed(12262,32), to_signed(12068,32), to_signed(69,32), to_signed(296,32), to_signed(55,32), to_signed(372,32), to_signed(11998,32), to_signed(2,32), to_signed(12218,32), to_signed(11974,32), to_signed(12282,32), to_signed(113,32), to_signed(12116,32), to_signed(318,32), to_signed(41,32), to_signed(241,32), to_signed(565,32), to_signed(12102,32), to_signed(12076,32), to_signed(12275,32), to_signed(14,32), to_signed(105,32), to_signed(21,32), to_signed(12249,32), to_signed(187,32), to_signed(11937,32), to_signed(12228,32), to_signed(107,32), to_signed(186,32), to_signed(12266,32), to_signed(11806,32), to_signed(12245,32), to_signed(47,32), to_signed(12199,32), to_signed(12227,32), to_signed(12288,32), to_signed(12175,32), to_signed(82,32), to_signed(11799,32), to_signed(12018,32), to_signed(206,32), to_signed(267,32), to_signed(74,32), to_signed(1,32), to_signed(71,32), to_signed(12232,32), to_signed(193,32), to_signed(12264,32), to_signed(11980,32), to_signed(12249,32), to_signed(12055,32), to_signed(12068,32), to_signed(373,32), to_signed(67,32), to_signed(111,32), to_signed(240,32), to_signed(171,32), to_signed(83,32), to_signed(12148,32), to_signed(136,32), to_signed(342,32), to_signed(88,32), to_signed(12276,32), to_signed(12257,32), to_signed(12183,32), to_signed(139,32), to_signed(12207,32), to_signed(12259,32), to_signed(467,32), to_signed(166,32), to_signed(85,32), to_signed(11851,32), to_signed(12005,32), to_signed(344,32), to_signed(12206,32), to_signed(170,32), to_signed(263,32), to_signed(11919,32), to_signed(12285,32), to_signed(24,32), to_signed(174,32), to_signed(12092,32), to_signed(11920,32), to_signed(11947,32), to_signed(12035,32), to_signed(12154,32), to_signed(89,32), to_signed(99,32), to_signed(165,32), to_signed(12222,32), to_signed(150,32), to_signed(544,32), to_signed(108,32));


  signal u : ram_type := (to_signed(13380, 32), to_signed(2111, 32), to_signed(4754, 32), to_signed(5327, 32), to_signed(10499, 32), to_signed(12902, 32), to_signed(8409, 32), to_signed(13827, 32), to_signed(20148, 32), to_signed(15176, 32), to_signed(4376, 32), to_signed(6918, 32), to_signed(10092, 32), to_signed(18881, 32), to_signed(20847, 32), to_signed(14802, 32), to_signed(1259, 32), to_signed(6283, 32), to_signed(996, 32), to_signed(16055, 32), to_signed(9280, 32), to_signed(3160, 32), to_signed(15542, 32), to_signed(21790, 32), to_signed(12603, 32), to_signed(19032, 32), to_signed(23889, 32), to_signed(14719, 32), to_signed(18006, 32), to_signed(10874, 32), to_signed(5797, 32), to_signed(1400, 32), to_signed(13631, 32), to_signed(2877, 32), to_signed(15866, 32), to_signed(18473, 32), to_signed(22534, 32), to_signed(19426, 32), to_signed(873, 32), to_signed(24332, 32), to_signed(17736, 32), to_signed(1088, 32), to_signed(2162, 32), to_signed(8822, 32), to_signed(18755, 32), to_signed(10304, 32), to_signed(24108, 32), to_signed(7552, 32), to_signed(6002, 32), to_signed(24485, 32), to_signed(14038, 32), to_signed(24274, 32), to_signed(3032, 32), to_signed(4881, 32), to_signed(979, 32), to_signed(24489, 32), to_signed(23230, 32), to_signed(11530, 32), to_signed(22636, 32), to_signed(941, 32), to_signed(8457, 32), to_signed(7829, 32), to_signed(13518, 32), to_signed(3864, 32), to_signed(19722, 32), to_signed(9337, 32), to_signed(22439, 32), to_signed(4030, 32), to_signed(14874, 32), to_signed(24026, 32), to_signed(9091, 32), to_signed(6638, 32), to_signed(19745, 32), to_signed(4002, 32), to_signed(5547, 32), to_signed(17267, 32), to_signed(12265, 32), to_signed(9220, 32), to_signed(23630, 32), to_signed(23952, 32), to_signed(24238, 32), to_signed(4526, 32), to_signed(1593, 32), to_signed(4808, 32), to_signed(4401, 32), to_signed(15633, 32), to_signed(7100, 32), to_signed(1196, 32), to_signed(19118, 32), to_signed(1451, 32), to_signed(7966, 32), to_signed(7754, 32), to_signed(15304, 32), to_signed(17765, 32), to_signed(11339, 32), to_signed(820, 32), to_signed(373, 32), to_signed(21646, 32), to_signed(18197, 32), to_signed(21325, 32), to_signed(10950, 32), to_signed(21940, 32), to_signed(11468, 32), to_signed(14604, 32), to_signed(22998, 32), to_signed(1988, 32), to_signed(6515, 32), to_signed(9001, 32), to_signed(8303, 32), to_signed(1915, 32), to_signed(9776, 32), to_signed(6917, 32), to_signed(12152, 32), to_signed(10321, 32), to_signed(19715, 32), to_signed(20867, 32), to_signed(9705, 32), to_signed(23172, 32), to_signed(7978, 32), to_signed(6833, 32), to_signed(392, 32), to_signed(17802, 32), to_signed(19533, 32), to_signed(23730, 32), to_signed(9191, 32), to_signed(9517, 32), to_signed(17075, 32), to_signed(10426, 32), to_signed(22390, 32), to_signed(9101, 32), to_signed(15107, 32), to_signed(1271, 32), to_signed(22739, 32), to_signed(1535, 32), to_signed(12520, 32), to_signed(14337, 32), to_signed(3857, 32), to_signed(2594, 32), to_signed(17734, 32), to_signed(18943, 32), to_signed(13846, 32), to_signed(10810, 32), to_signed(2447, 32), to_signed(12722, 32), to_signed(12300, 32), to_signed(20352, 32), to_signed(17120, 32), to_signed(18727, 32), to_signed(18476, 32), to_signed(2683, 32), to_signed(1505, 32), to_signed(10004, 32), to_signed(20018, 32), to_signed(5355, 32), to_signed(21733, 32), to_signed(19062, 32), to_signed(9304, 32), to_signed(9900, 32), to_signed(18281, 32), to_signed(7541, 32), to_signed(9398, 32), to_signed(18552, 32), to_signed(1425, 32), to_signed(15990, 32), to_signed(13773, 32), to_signed(15149, 32), to_signed(8104, 32), to_signed(5991, 32), to_signed(19278, 32), to_signed(5552, 32), to_signed(6848, 32), to_signed(10259, 32), to_signed(22547, 32), to_signed(23809, 32), to_signed(10443, 32), to_signed(1977, 32), to_signed(674, 32), to_signed(22754, 32), to_signed(14181, 32), to_signed(10617, 32), to_signed(10880, 32), to_signed(11449, 32), to_signed(19849, 32), to_signed(2830, 32), to_signed(13908, 32), to_signed(18198, 32), to_signed(21469, 32), to_signed(13983, 32), to_signed(2025, 32), to_signed(16059, 32), to_signed(13701, 32), to_signed(4250, 32), to_signed(24061, 32), to_signed(905, 32), to_signed(1358, 32), to_signed(10118, 32), to_signed(19154, 32), to_signed(8550, 32), to_signed(4200, 32), to_signed(23230, 32), to_signed(14346, 32), to_signed(554, 32), to_signed(855, 32), to_signed(5617, 32), to_signed(701, 32), to_signed(15431, 32), to_signed(6966, 32), to_signed(16578, 32), to_signed(14057, 32), to_signed(3785, 32), to_signed(2766, 32), to_signed(3544, 32), to_signed(14476, 32), to_signed(10612, 32), to_signed(129, 32), to_signed(16888, 32), to_signed(15911, 32), to_signed(1546, 32), to_signed(6703, 32), to_signed(17307, 32), to_signed(10114, 32), to_signed(20350, 32), to_signed(11216, 32), to_signed(10667, 32), to_signed(17946, 32), to_signed(12007, 32), to_signed(15387, 32), to_signed(206, 32), to_signed(9538, 32), to_signed(1339, 32), to_signed(8146, 32), to_signed(17423, 32), to_signed(2617, 32), to_signed(9883, 32), to_signed(21079, 32), to_signed(18508, 32), to_signed(8847, 32), to_signed(150, 32), to_signed(20876, 32), to_signed(23964, 32), to_signed(20150, 32), to_signed(13533, 32), to_signed(18288, 32), to_signed(12926, 32), to_signed(19381, 32), to_signed(9946, 32), to_signed(4064, 32), to_signed(12553, 32), to_signed(2078, 32), to_signed(8331, 32), to_signed(7634, 32), to_signed(18978, 32), to_signed(9864, 32), to_signed(8763, 32), to_signed(14147, 32), to_signed(7190, 32), to_signed(19008, 32), to_signed(7157, 32), to_signed(13285, 32), to_signed(10151, 32), to_signed(7649, 32), to_signed(11493, 32), to_signed(3061, 32), to_signed(9322, 32), to_signed(15970, 32), to_signed(3593, 32), to_signed(9858, 32), to_signed(7873, 32), to_signed(11055, 32), to_signed(20532, 32), to_signed(14999, 32), to_signed(19809, 32), to_signed(14741, 32), to_signed(2216, 32), to_signed(3919, 32), to_signed(15006, 32), to_signed(17844, 32), to_signed(24474, 32), to_signed(22993, 32), to_signed(20853, 32), to_signed(10504, 32), to_signed(24527, 32), to_signed(21515, 32), to_signed(16082, 32), to_signed(11774, 32), to_signed(8941, 32), to_signed(11829, 32), to_signed(24010, 32), to_signed(10178, 32), to_signed(22316, 32), to_signed(17426, 32), to_signed(3448, 32), to_signed(11618, 32), to_signed(20185, 32), to_signed(7217, 32), to_signed(11844, 32), to_signed(3095, 32), to_signed(20948, 32), to_signed(323, 32), to_signed(7078, 32), to_signed(3097, 32), to_signed(9811, 32), to_signed(16190, 32), to_signed(24486, 32), to_signed(2235, 32), to_signed(9252, 32), to_signed(14981, 32), to_signed(2652, 32), to_signed(12844, 32), to_signed(23088, 32), to_signed(12529, 32), to_signed(18786, 32), to_signed(19283, 32), to_signed(11486, 32), to_signed(6213, 32), to_signed(18721, 32), to_signed(24376, 32), to_signed(19953, 32), to_signed(17593, 32), to_signed(21636, 32), to_signed(1406, 32), to_signed(4421, 32), to_signed(6328, 32), to_signed(18026, 32), to_signed(10302, 32), to_signed(1630, 32), to_signed(1253, 32), to_signed(11792, 32), to_signed(12976, 32), to_signed(12789, 32), to_signed(24545, 32), to_signed(18225, 32), to_signed(20007, 32), to_signed(18784, 32), to_signed(4693, 32), to_signed(16583, 32), to_signed(15521, 32), to_signed(11056, 32), to_signed(16277, 32), to_signed(9533, 32), to_signed(20500, 32), to_signed(15975, 32), to_signed(20234, 32), to_signed(5904, 32), to_signed(844, 32), to_signed(21255, 32), to_signed(9833, 32), to_signed(21899, 32), to_signed(3051, 32), to_signed(17220, 32), to_signed(4728, 32), to_signed(15495, 32), to_signed(15489, 32), to_signed(8801, 32), to_signed(5349, 32), to_signed(11263, 32), to_signed(17823, 32), to_signed(24057, 32), to_signed(830, 32), to_signed(19981, 32), to_signed(1139, 32), to_signed(10986, 32), to_signed(18656, 32), to_signed(7757, 32), to_signed(6930, 32), to_signed(23615, 32), to_signed(5727, 32), to_signed(15304, 32), to_signed(9441, 32), to_signed(6888, 32), to_signed(21698, 32), to_signed(21095, 32), to_signed(20557, 32), to_signed(5824, 32), to_signed(5371, 32), to_signed(4927, 32), to_signed(16052, 32), to_signed(11454, 32), to_signed(2979, 32), to_signed(20655, 32), to_signed(5465, 32), to_signed(8272, 32), to_signed(8566, 32), to_signed(20057, 32), to_signed(16983, 32), to_signed(18721, 32), to_signed(9545, 32), to_signed(4968, 32), to_signed(10437, 32), to_signed(8364, 32), to_signed(3228, 32), to_signed(24545, 32), to_signed(17615, 32), to_signed(13391, 32), to_signed(11267, 32), to_signed(10077, 32), to_signed(6489, 32), to_signed(19736, 32), to_signed(14430, 32), to_signed(14898, 32), to_signed(23672, 32), to_signed(2255, 32), to_signed(6622, 32), to_signed(3300, 32), to_signed(4034, 32), to_signed(941, 32), to_signed(18918, 32), to_signed(4776, 32), to_signed(15247, 32), to_signed(23234, 32), to_signed(10075, 32), to_signed(12161, 32), to_signed(13921, 32), to_signed(23788, 32), to_signed(22592, 32), to_signed(4419, 32), to_signed(24344, 32), to_signed(15374, 32), to_signed(1656, 32), to_signed(6963, 32), to_signed(10857, 32), to_signed(21531, 32), to_signed(1454, 32), to_signed(1139, 32), to_signed(8398, 32), to_signed(20501, 32), to_signed(6888, 32), to_signed(9117, 32), to_signed(7065, 32), to_signed(14835, 32), to_signed(15259, 32), to_signed(1087, 32), to_signed(13888, 32), to_signed(18095, 32), to_signed(2325, 32), to_signed(3105, 32), to_signed(563, 32), to_signed(6637, 32), to_signed(6228, 32), to_signed(402, 32), to_signed(12109, 32), to_signed(3383, 32), to_signed(24568, 32), to_signed(12969, 32), to_signed(842, 32), to_signed(9051, 32), to_signed(16691, 32), to_signed(3750, 32), to_signed(13897, 32), to_signed(4639, 32), to_signed(19452, 32), to_signed(24409, 32), to_signed(20228, 32), to_signed(2860, 32), to_signed(22037, 32), to_signed(17366, 32), to_signed(13136, 32), to_signed(13600, 32), to_signed(4209, 32), to_signed(7554, 32), to_signed(18843, 32), to_signed(23132, 32), to_signed(7681, 32), to_signed(17063, 32), to_signed(18781, 32), to_signed(21131, 32), to_signed(24117, 32), to_signed(14563, 32), to_signed(17848, 32), to_signed(10324, 32), to_signed(13657, 32), to_signed(9509, 32), to_signed(5443, 32), to_signed(6959, 32), to_signed(2042, 32), to_signed(24541, 32), to_signed(1117, 32), to_signed(20949, 32), to_signed(16314, 32), to_signed(17810, 32), to_signed(4644, 32), to_signed(24375, 32), to_signed(7482, 32), to_signed(10078, 32), to_signed(14121, 32), to_signed(12824, 32), to_signed(16666, 32), to_signed(13193, 32), to_signed(23090, 32), to_signed(21169, 32), to_signed(21380, 32), to_signed(7352, 32), to_signed(3072, 32), to_signed(1569, 32), to_signed(4134, 32), to_signed(18197, 32), to_signed(14774, 32), to_signed(19088, 32), to_signed(15124, 32), to_signed(8294, 32), to_signed(10517, 32), to_signed(5715, 32), to_signed(24510, 32), to_signed(6698, 32), to_signed(23611, 32), to_signed(1451, 32), to_signed(15999, 32), to_signed(11675, 32), to_signed(18479, 32), to_signed(14586, 32), to_signed(15192, 32), to_signed(1314, 32));


  signal sc1 : ram_type := (to_signed(3, 32), to_signed(-5, 32), to_signed(3, 32), to_signed(-4, 32), to_signed(3, 32), to_signed(2, 32), to_signed(3, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(3, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(3, 32), to_signed(5, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(4, 32), to_signed(2, 32), to_signed(1, 32), to_signed(1, 32), to_signed(3, 32), to_signed(4, 32), to_signed(1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(3, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(1, 32), to_signed(3, 32), to_signed(3, 32), to_signed(-5, 32), to_signed(-1, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(2, 32), to_signed(2, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(3, 32), to_signed(4, 32), to_signed(2, 32), to_signed(2, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-4, 32), to_signed(-5, 32), to_signed(6, 32), to_signed(2, 32), to_signed(5, 32), to_signed(2, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(1, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(3, 32), to_signed(3, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(4, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-6, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-5, 32), to_signed(3, 32), to_signed(2, 32), to_signed(1, 32), to_signed(2, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(3, 32), to_signed(-6, 32), to_signed(1, 32), to_signed(0, 32), to_signed(1, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(4, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(2, 32), to_signed(3, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-5, 32), to_signed(3, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(-1, 32), to_signed(6, 32), to_signed(7, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(0, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(3, 32), to_signed(2, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(0, 32), to_signed(0, 32), to_signed(2, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(0, 32), to_signed(1, 32), to_signed(4, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(6, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(0, 32), to_signed(2, 32), to_signed(1, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(-4, 32), to_signed(-5, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(1, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-6, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(0, 32), to_signed(5, 32), to_signed(5, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(3, 32), to_signed(3, 32), to_signed(0, 32), to_signed(-7, 32), to_signed(3, 32), to_signed(1, 32), to_signed(2, 32), to_signed(3, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(3, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(4, 32), to_signed(5, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(-8, 32), to_signed(-1, 32), to_signed(4, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(4, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(3, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(5, 32), to_signed(-1, 32), to_signed(3, 32), to_signed(4, 32), to_signed(-1, 32), to_signed(3, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(3, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-5, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(0, 32), to_signed(3, 32), to_signed(4, 32), to_signed(1, 32), to_signed(5, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(3, 32), to_signed(1, 32), to_signed(3, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(2, 32), to_signed(2, 32), to_signed(3, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-3, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-3, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-4, 32), to_signed(-3, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-5, 32), to_signed(4, 32), to_signed(3, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-5, 32), to_signed(2, 32), to_signed(-7, 32), to_signed(-1, 32), to_signed(0, 32), to_signed(0, 32), to_signed(3, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(3, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(-3, 32), to_signed(0, 32), to_signed(-5, 32), to_signed(-5, 32), to_signed(1, 32), to_signed(-1, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(2, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(0, 32), to_signed(0, 32), to_signed(3, 32), to_signed(1, 32), to_signed(0, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(3, 32), to_signed(-4, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-3, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(1, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(-1, 32), to_signed(-3, 32));


  signal sc2 : ram_type := (to_signed(6, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(6, 32), to_signed(8, 32), to_signed(12, 32), to_signed(-4, 32), to_signed(8, 32), to_signed(6, 32), to_signed(-6, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(4, 32), to_signed(0, 32), to_signed(8, 32), to_signed(4, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(8, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(0, 32), to_signed(14, 32), to_signed(-8, 32), to_signed(10, 32), to_signed(2, 32), to_signed(10, 32), to_signed(2, 32), to_signed(2, 32), to_signed(4, 32), to_signed(10, 32), to_signed(2, 32), to_signed(6, 32), to_signed(-2, 32), to_signed(-8, 32), to_signed(16, 32), to_signed(2, 32), to_signed(-8, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(16, 32), to_signed(2, 32), to_signed(-14, 32), to_signed(14, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(2, 32), to_signed(0, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-1, 32), to_signed(8, 32), to_signed(6, 32), to_signed(4, 32), to_signed(-8, 32), to_signed(-6, 32), to_signed(10, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(1, 32), to_signed(4, 32), to_signed(6, 32), to_signed(4, 32), to_signed(2, 32), to_signed(4, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(-8, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(10, 32), to_signed(4, 32), to_signed(2, 32), to_signed(4, 32), to_signed(4, 32), to_signed(0, 32), to_signed(8, 32), to_signed(2, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(14, 32), to_signed(5, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(2, 32), to_signed(10, 32), to_signed(12, 32), to_signed(-4, 32), to_signed(6, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(8, 32), to_signed(-6, 32), to_signed(8, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(2, 32), to_signed(4, 32), to_signed(8, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(2, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(13, 32), to_signed(0, 32), to_signed(6, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(8, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-7, 32), to_signed(6, 32), to_signed(4, 32), to_signed(8, 32), to_signed(2, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(-8, 32), to_signed(-4, 32), to_signed(8, 32), to_signed(-2, 32), to_signed(12, 32), to_signed(8, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(2, 32), to_signed(0, 32), to_signed(6, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(2, 32), to_signed(1, 32), to_signed(2, 32), to_signed(0, 32), to_signed(4, 32), to_signed(2, 32), to_signed(6, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(8, 32), to_signed(4, 32), to_signed(6, 32), to_signed(8, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-6, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(2, 32), to_signed(10, 32), to_signed(9, 32), to_signed(-2, 32), to_signed(-8, 32), to_signed(12, 32), to_signed(6, 32), to_signed(0, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(0, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(4, 32), to_signed(2, 32), to_signed(8, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(0, 32), to_signed(6, 32), to_signed(2, 32), to_signed(2, 32), to_signed(4, 32), to_signed(8, 32), to_signed(-6, 32), to_signed(0, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(9, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(4, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(10, 32), to_signed(6, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(10, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(10, 32), to_signed(-6, 32), to_signed(1, 32), to_signed(2, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(1, 32), to_signed(-4, 32), to_signed(12, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(2, 32), to_signed(2, 32), to_signed(-1, 32), to_signed(4, 32), to_signed(0, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-6, 32), to_signed(8, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(4, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(-8, 32), to_signed(6, 32), to_signed(2, 32), to_signed(1, 32), to_signed(6, 32), to_signed(-5, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(6, 32), to_signed(2, 32), to_signed(8, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(2, 32), to_signed(2, 32), to_signed(2, 32), to_signed(10, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-6, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(-12, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(-10, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(-6, 32), to_signed(-6, 32), to_signed(8, 32), to_signed(-2, 32), to_signed(-6, 32), to_signed(12, 32), to_signed(-14, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(2, 32), to_signed(-7, 32), to_signed(6, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-2, 32), to_signed(10, 32), to_signed(1, 32), to_signed(2, 32), to_signed(4, 32), to_signed(-8, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-10, 32), to_signed(-8, 32), to_signed(7, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(10, 32), to_signed(-16, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(2, 32), to_signed(-12, 32), to_signed(-2, 32), to_signed(8, 32), to_signed(6, 32), to_signed(-2, 32), to_signed(4, 32), to_signed(2, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(8, 32), to_signed(-8, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-9, 32), to_signed(-4, 32), to_signed(4, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(-14, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(2, 32), to_signed(0, 32), to_signed(6, 32), to_signed(12, 32), to_signed(4, 32), to_signed(0, 32), to_signed(-12, 32), to_signed(-12, 32), to_signed(2, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(6, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(-10, 32), to_signed(-2, 32), to_signed(-8, 32), to_signed(-14, 32), to_signed(4, 32), to_signed(-10, 32), to_signed(4, 32), to_signed(-10, 32), to_signed(-4, 32), to_signed(6, 32), to_signed(-10, 32), to_signed(2, 32), to_signed(-12, 32), to_signed(2, 32), to_signed(-8, 32), to_signed(10, 32), to_signed(-10, 32), to_signed(0, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(-10, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(1, 32), to_signed(0, 32), to_signed(4, 32), to_signed(-4, 32), to_signed(8, 32), to_signed(-4, 32), to_signed(-6, 32), to_signed(0, 32), to_signed(-6, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(2, 32), to_signed(-8, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(-8, 32), to_signed(4, 32), to_signed(-6, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(-6, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(-10, 32), to_signed(-4, 32), to_signed(-6, 32), to_signed(10, 32), to_signed(-5, 32), to_signed(2, 32), to_signed(-4, 32), to_signed(14, 32), to_signed(-6, 32), to_signed(4, 32), to_signed(-8, 32), to_signed(-10, 32), to_signed(8, 32), to_signed(1, 32), to_signed(-2, 32), to_signed(-8, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-6, 32), to_signed(-9, 32), to_signed(2, 32), to_signed(-6, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(6, 32), to_signed(0, 32), to_signed(-14, 32), to_signed(-4, 32), to_signed(12, 32), to_signed(-2, 32), to_signed(-6, 32), to_signed(0, 32), to_signed(0, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-4, 32), to_signed(-8, 32), to_signed(-10, 32), to_signed(2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(-2, 32), to_signed(-2, 32), to_signed(0, 32), to_signed(2, 32), to_signed(6, 32), to_signed(0, 32), to_signed(-4, 32), to_signed(-18, 32), to_signed(-4, 32), to_signed(-2, 32), to_signed(-4, 32), to_signed(-8, 32), to_signed(-2, 32));


  signal reset           : std_logic;
  signal rejection       : std_logic;
  signal coeff_sc_addr   : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0) := (others => '0');
  signal coeff_sc1       : std_logic_vector(MAX_RES_WIDTH-1 downto 0)                         := (others => '0');
  signal coeff_sc1_valid : std_logic                                                          := '0';
  signal coeff_sc2       : std_logic_vector(MAX_RES_WIDTH-1 downto 0)                         := (others => '0');
  signal coeff_sc2_valid : std_logic                                                          := '0';
  signal delay_temp_ram  : integer range 0 to 63                                              := 10;
  signal u_data          : std_logic_vector(PRIME_P'length+1-1 downto 0)                      := (others => '0');
  signal u_addr          : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0) := (others => '0');
  signal y1_data         : std_logic_vector(PRIME_P'length-1 downto 0)                        := (others => '0');
  signal y1_addr         : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0) := (others => '0');
  signal y2_data         : std_logic_vector(PRIME_P'length-1 downto 0)                        := (others => '0');
  signal y2_addr         : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0) := (others => '0');
  signal z2_final        : std_logic_vector(1 downto 0)                                       := (others => '0');
  signal z2_final_addr   : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0)           := (others => '0');
  signal z2_final_valid  : std_logic                                                          := '0';

  signal z1_final        : std_logic_vector(PRIME_P'length-1 downto 0)                                       := (others => '0');
  signal z1_final_addr   : std_logic_vector(integer(ceil(log2(real(N_ELEMENTS))))-1 downto 0)           := (others => '0');
  signal z1_final_valid  : std_logic                                                          := '0';
begin

  process (clk)
  begin  -- process
    if rising_edge(clk) then
      
      u_data  <= std_logic_vector(resize(unsigned(u(to_integer(unsigned(u_addr)))),u_data'length));
      y1_data <= std_logic_vector(resize(unsigned(y1(to_integer(unsigned(y1_addr)))),y1_data'length));
      y2_data <= std_logic_vector(resize(unsigned(y2(to_integer(unsigned(y2_addr)))),y2_data'length));
      
    end if;
  end process;


  rejection_module_1 : entity work.rejection_module
    generic map (
      N_ELEMENTS             => N_ELEMENTS,
      PRIME_P_WIDTH          => PRIME_P_WIDTH,
      PRIME_P                => PRIME_P,
      ZETA                   => ZETA,
      D_BLISS                => D_BLISS,
      MODULUS_P_BLISS        => MODULUS_P_BLISS,
      MAX_RES_WIDTH_COEFF_SC => MAX_RES_WIDTH,
      CORES                  => CORES,
      KAPPA                  => KAPPA,
      WIDTH_S1               => WIDTH_S1,
      WIDTH_S2               => WIDTH_S2,
      INIT_TABLE             => INIT_TABLE,
      c_delay                => c_delay,
      MAX_RES_WIDTH          => MAX_RES_WIDTH
      )
    port map (
      clk             => clk,
      reset           => reset,
      rejection       => rejection,
      coeff_sc_addr   => coeff_sc_addr,
      coeff_sc1       => coeff_sc1,
      coeff_sc1_valid => coeff_sc1_valid,
      coeff_sc2       => coeff_sc2,
      coeff_sc2_valid => coeff_sc2_valid,
      delay_temp_ram  => delay_temp_ram,
      u_data          => u_data,
      u_addr          => u_addr,
      y1_data         => y1_data,
      y1_addr         => y1_addr,
      y2_data         => y2_data,
      y2_addr         => y2_addr,
      z1_final        => z1_final,
      z1_final_addr   => z1_final_addr,
      z1_final_valid  => z1_final_valid,
      z2_final        => z2_final,
      z2_final_addr   => z2_final_addr,
      z2_final_valid  => z2_final_valid
      );

  
  clk_process : process
  begin
    if end_of_simulation = '0' then
      clk           <= '0';
      wait for clk_period/2;
      clk           <= '1';
      wait for clk_period/2;
      cycle_counter <= cycle_counter+1;
    end if;
  end process;
  end_of_simulation_out <= end_of_simulation;



  -- Stimulus process
  stim_proc : process
  begin
    -- hold reset state for 100 ns.
    wait for 100 ns;


    for i in 0 to 511 loop
      coeff_sc_addr <=std_logic_vector( to_unsigned(i,coeff_sc_addr'length));
      coeff_sc1_valid <= '1';
      coeff_sc1       <= std_logic_vector(resize(unsigned(sc1(i)), coeff_sc1'length));
      coeff_sc2_valid <= '1';
      coeff_sc2       <= std_logic_vector(resize(unsigned(sc2(i)), coeff_sc2'length));
      wait for clk_period;
    end loop;  -- i 
    coeff_sc2_valid <= '0';
    coeff_sc1_valid <= '0';

    wait for clk_period*1000;


    if error_happened = '1' then
      report "ERROR";
    else
      report "OK";
    end if;

    end_of_simulation <= '1';
    wait;

    -- insert stimulus here 

    wait;
  end process;




  
end;
