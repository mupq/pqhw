--/****************************************************************************/
--Copyright (C) by Thomas P�ppelmann and the Hardware Security Group of Ruhr-Universitaet Bochum. 
--All rights reserved.
--This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. 
--Please see licence.rtf and readme.txt for licence and further instructions.
--/****************************************************************************/

--
--      Package File Template
--
--      Purpose: This package defines supplemental types, subtypes, 
--               constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;



package cdt_sampler_pkg is

  constant MAX_REVERSE_ENTRY : integer := 400;

  type reverse_entry_type is array (0 to 1) of integer range 0 to MAX_REVERSE_ENTRY;
  type reverse_table_type is array (natural range <>) of reverse_entry_type;

  constant NUM_INTERVALS : integer := 16;
  constant MAX_INTERVAL  : integer := 4000;
  type     intervals_type is array (0 to NUM_INTERVALS-1) of integer range 0 to MAX_INTERVAL;
  type     max_tables_type is array (0 to NUM_INTERVALS-1) of integer range 0 to MAX_INTERVAL;


  subtype exp_array_entry is integer range 0 to 192;
  type    exp_array_type is array (natural range <>) of exp_array_entry;





  function get_cdt_max_index (param      : integer) return integer;
  function get_cdt_max_byte (param       : integer) return integer;
  function get_cdt_max_byte_table (param : integer) return integer;
  function get_reverse_table(param       : integer) return reverse_table_type;
  function get_get_mul_factor(param      : integer) return integer;
  function get_intervals_table(param     : integer) return intervals_type;
  function get_intervals_table_max(param : integer) return intervals_type;
  function get_max_ram (param            : integer) return integer;
  function get_sigma(param               : integer) return real;
  function get_max_sigma(param           : integer) return integer;
  function get_gauss_prob(x, sigma       : real) return real;
  function get_absolute(x                : real) return real;
  function get_exponent_table(param      : integer) return exp_array_type;

  function get_max_exponent(param : integer) return integer;

  
end cdt_sampler_pkg;

package body cdt_sampler_pkg is

  function get_sigma(param : integer) return real is
  begin
    if param = 1 then
      return 215.7277372731568368513;
    elsif param = 3 then
      return 250.5499310849656176028;
    elsif param = 4 then
      return 270.9336542918780746282;
    end if;
  end get_sigma;


  function get_max_sigma(param : integer) return integer is
  begin
    return get_cdt_max_index(param)+get_get_mul_factor(param)*get_cdt_max_index(param);
  end get_max_sigma;


  function get_get_mul_factor(param : integer) return integer is
  begin
    if param = 1 then
      return 11;
    elsif param = 3 then
      return 12;
    elsif param = 4 then
      return 11;
    end if;
  end get_get_mul_factor;


  function get_cdt_max_byte_table (param : integer) return integer is
  begin
    if param = 1 then
      return 8;
    elsif param = 3 then
      return 10;
    elsif param = 4 then
      return 13;
    end if;
  end get_cdt_max_byte_table;


  function get_cdt_max_byte (param : integer) return integer is
  begin
    if param = 1 then
      return 35;
    elsif param = 3 then
      return 35;
    elsif param = 4 then
      return 35;
    end if;
  end get_cdt_max_byte;


  function get_intervals_table_max(param : integer) return intervals_type is
    constant max_table_1 : intervals_type := (262, 262, 235, 223, 202, 180, 157, 125, 86, 0, 0, 0, 0, 0, 0, 0);
    constant max_table_3 : intervals_type := (371, 308, 292, 279, 259, 236, 215, 192, 167, 121, 94, 0, 0, 0, 0, 0);
    constant max_table_4 : intervals_type := (400, 393, 383, 364, 344, 332, 302, 278, 246, 226, 197, 155, 111, 0, 0, 0);

  begin
    if param = 1 then
      return max_table_1;
    end if;
    if param = 3 then
      return max_table_3;
    elsif param = 4 then
      return max_table_4;
    end if;
  end get_intervals_table_max;



  function get_reverse_table(param : integer) return reverse_table_type is
    constant reverse_table_bliss_1 : reverse_table_type := ((56, 262), (52, 57), (49, 53), (47, 50), (46, 48), (44, 47), (43, 45), (42, 44), (41, 43), (40, 42), (40, 41), (39, 41), (38, 40), (38, 39), (37, 39), (36, 38), (36, 37), (35, 37), (35, 36), (34, 36), (34, 35), (34, 35), (33, 35), (33, 34), (32, 34), (32, 33), (32, 33), (31, 33), (31, 32), (31, 32), (30, 32), (30, 31), (30, 31), (29, 31), (29, 30), (29, 30), (28, 30), (28, 29), (28, 29), (28, 29), (27, 29), (27, 28), (27, 28), (27, 28), (26, 28), (26, 27), (26, 27), (26, 27), (26, 27), (25, 27), (25, 26), (25, 26), (25, 26), (24, 26), (24, 25), (24, 25), (24, 25), (24, 25), (23, 25), (23, 24), (23, 24), (23, 24), (23, 24), (22, 24), (22, 23), (22, 23), (22, 23), (22, 23), (22, 23), (21, 23), (21, 22), (21, 22), (21, 22), (21, 22), (21, 22), (20, 22), (20, 21), (20, 21), (20, 21), (20, 21), (20, 21), (19, 21), (19, 20), (19, 20), (19, 20), (19, 20), (19, 20), (18, 20), (18, 19), (18, 19), (18, 19), (18, 19), (18, 19), (18, 19), (17, 19), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (16, 18), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (15, 17), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (14, 16), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (13, 15), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (12, 14), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (11, 13), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (10, 12), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (9, 11), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (8, 10), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (7, 9), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (6, 8), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (5, 7), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (4, 6), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (3, 5), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (2, 4), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (1, 3), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (0, 2), (0, 1), (0, 1), (0, 1), (0, 1), (0, 1));

    constant reverse_table_bliss_3 : reverse_table_type := ((60, 317), (55, 61), (52, 56), (50, 53), (49, 51), (47, 50), (46, 48), (45, 47), (44, 46), (43, 45), (42, 44), (41, 43), (41, 42), (40, 42), (39, 41), (39, 40), (38, 40), (38, 39), (37, 39), (37, 38), (36, 38), (36, 37), (35, 37), (35, 36), (34, 36), (34, 35), (34, 35), (33, 35), (33, 34), (33, 34), (32, 34), (32, 33), (32, 33), (31, 33), (31, 32), (31, 32), (30, 32), (30, 31), (30, 31), (29, 31), (29, 30), (29, 30), (29, 30), (28, 30), (28, 29), (28, 29), (28, 29), (27, 29), (27, 28), (27, 28), (27, 28), (26, 28), (26, 27), (26, 27), (26, 27), (26, 27), (25, 27), (25, 26), (25, 26), (25, 26), (25, 26), (24, 26), (24, 25), (24, 25), (24, 25), (24, 25), (23, 25), (23, 24), (23, 24), (23, 24), (23, 24), (22, 24), (22, 23), (22, 23), (22, 23), (22, 23), (22, 23), (21, 23), (21, 22), (21, 22), (21, 22), (21, 22), (21, 22), (20, 22), (20, 21), (20, 21), (20, 21), (20, 21), (20, 21), (19, 21), (19, 20), (19, 20), (19, 20), (19, 20), (19, 20), (18, 20), (18, 19), (18, 19), (18, 19), (18, 19), (18, 19), (18, 19), (17, 19), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (16, 18), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (15, 17), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (14, 16), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (13, 15), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (12, 14), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (11, 13), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (10, 12), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (9, 11), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (8, 10), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (7, 9), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (6, 8), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (5, 7), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (4, 6), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (3, 5), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (2, 4), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (1, 3), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (0, 2), (0, 1), (0, 1), (0, 1), (0, 1));

    constant reverse_table_bliss_4 : reverse_table_type := ((71, 400), (65, 72), (62, 66), (59, 63), (57, 60), (56, 58), (54, 57), (53, 55), (52, 54), (51, 53), (50, 52), (49, 51), (48, 50), (47, 49), (46, 48), (46, 47), (45, 47), (44, 46), (44, 45), (43, 45), (43, 44), (42, 44), (42, 43), (41, 43), (41, 42), (40, 42), (40, 41), (39, 41), (39, 40), (38, 40), (38, 39), (38, 39), (37, 39), (37, 38), (36, 38), (36, 37), (36, 37), (35, 37), (35, 36), (35, 36), (34, 36), (34, 35), (34, 35), (34, 35), (33, 35), (33, 34), (33, 34), (32, 34), (32, 33), (32, 33), (31, 33), (31, 32), (31, 32), (31, 32), (30, 32), (30, 31), (30, 31), (30, 31), (29, 31), (29, 30), (29, 30), (29, 30), (28, 30), (28, 29), (28, 29), (28, 29), (28, 29), (27, 29), (27, 28), (27, 28), (27, 28), (26, 28), (26, 27), (26, 27), (26, 27), (26, 27), (25, 27), (25, 26), (25, 26), (25, 26), (25, 26), (24, 26), (24, 25), (24, 25), (24, 25), (24, 25), (23, 25), (23, 24), (23, 24), (23, 24), (23, 24), (22, 24), (22, 23), (22, 23), (22, 23), (22, 23), (22, 23), (21, 23), (21, 22), (21, 22), (21, 22), (21, 22), (21, 22), (20, 22), (20, 21), (20, 21), (20, 21), (20, 21), (20, 21), (19, 21), (19, 20), (19, 20), (19, 20), (19, 20), (19, 20), (18, 20), (18, 19), (18, 19), (18, 19), (18, 19), (18, 19), (17, 19), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (17, 18), (16, 18), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (16, 17), (15, 17), (15, 16), (15, 16), (15, 16), (15, 16), (15, 16), (14, 16), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (14, 15), (13, 15), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (13, 14), (12, 14), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (12, 13), (11, 13), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (11, 12), (10, 12), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (10, 11), (9, 11), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (9, 10), (8, 10), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (8, 9), (7, 9), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (7, 8), (6, 8), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (6, 7), (5, 7), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (5, 6), (4, 6), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (4, 5), (3, 5), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (3, 4), (2, 4), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (2, 3), (1, 3), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (1, 2), (0, 2), (0, 1), (0, 1), (0, 1), (0, 1));
    
  begin
    if param = 1 then
      return reverse_table_bliss_1;
    elsif param = 3 then
      return reverse_table_bliss_3;
    elsif param = 4 then
      return reverse_table_bliss_4;
    end if;
  end get_reverse_table;





  function get_exponent_table(param : integer) return exp_array_type is
    
    constant exp_array_1 : exp_array_type := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 , 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16);

    constant exp_array_3_no_divided : exp_array_type := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 112, 112, 112, 112, 112, 112, 112, 112, 112, 120, 120, 120, 120, 120, 120, 120, 120, 120, 128, 128, 128, 128, 128, 128, 128, 128, 136, 136, 136, 136, 136, 136, 136, 136, 136, 144, 144, 144, 144, 144, 144, 144, 144, 152, 152, 152, 152, 152, 152, 152, 152, 160, 160, 160, 160, 160, 160, 160, 168, 168, 168);

    variable exp_array_3 : exp_array_type(0 to exp_array_3_no_divided'length-1);

    constant exp_array_4_no_divided : exp_array_type := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 144, 144, 144, 144, 144, 144, 144, 144, 144, 152, 152, 152, 152, 152, 152, 152, 152, 152, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 168, 168, 168, 168, 168, 168, 168, 168, 176, 176, 176, 176, 176, 176, 176, 176, 176, 184, 184, 184, 184, 184, 184, 184, 184, 184, 192, 192, 192);

    variable exp_array_4 : exp_array_type(0 to exp_array_4_no_divided'length-1);
    
  begin
    if param = 1 then
      return exp_array_1;
    elsif param = 3 then
      for i in exp_array_3_no_divided'range loop
        exp_array_3(i) := exp_array_3_no_divided(i)/8;
      end loop;  -- i
      return exp_array_3;
    elsif param = 4 then
      for i in exp_array_4_no_divided'range loop
        exp_array_4(i) := exp_array_4_no_divided(i)/8;
      end loop;  -- i
      return exp_array_4;
    end if;
  end get_exponent_table;


  -----------------------------------------------------------------------------
  -- Parameter independent part
  -----------------------------------------------------------------------------
  function get_max_exponent (param : integer) return integer is
    constant exp_array : exp_array_type :=  get_exponent_table(param);
  begin
    return exp_array(exp_array'length-1);
  end;


  function get_max_ram (param : integer) return integer is
    variable max_table : intervals_type;
    variable val       : integer := 0;
  begin
    max_table := get_intervals_table_max(param);
    val       := 0;                     --Exponents
    for i in 0 to intervals_type'right loop
      val := val + max_table(i);
    end loop;

    return val;
  end get_max_ram;


  function get_intervals_table(param : integer) return intervals_type is
    variable intervals : intervals_type;
    variable max_table : intervals_type;
  begin

    --Get the max table
    max_table    := get_intervals_table_max(param);
    intervals(0) := 0;                  --Exponents
    for i in 0 to intervals_type'right-1 loop
      if max_table(i) /= 0 then
        intervals(i+1) := intervals(i)+max_table(i);
      else
        intervals(i+1) := 0;
      end if;
    end loop;  -- i

    return intervals;
  end get_intervals_table;



  function get_cdt_max_index (param : integer) return integer is
    variable max_table : intervals_type;
  begin
    max_table := get_intervals_table_max(param);
    return max_table(0);
  end get_cdt_max_index;



  function get_absolute(x : real) return real is
  begin
    if x < 0.0 then
      return -x;
    end if;

    return x;
  end get_absolute;

  function get_gauss_prob(x, sigma : real) return real is
    variable divisor  : real := 0.0;
    variable dividend : real := 0.0;
    variable exponent : real := 0.0;
  begin
    divisor  := SQRT(2.0*MATH_PI)*sigma;
    exponent := -x*x/(2.0*sigma*sigma);
    dividend := MATH_E**(exponent);
    return dividend/divisor;
  end get_gauss_prob;




  
end cdt_sampler_pkg;






















-------------------------------------------------------------------------------
-- 
-------------------------------------------------------------------------------
--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--use ieee.numeric_std.all;


--package cdt_sampler_pkg is

--  type reverse_entry_type is array (0 to 1) of integer;
--  type reverse_table_type is array (0 to 255) of unsigned(15 downto 0);

--  constant NUM_INTERVALS : integer := 16;
--  constant MAX_INTERVAL  : integer := 2314;
--  type     intervals_type is array (0 to NUM_INTERVALS-1) of integer;
--  type     max_tables_type is array (0 to NUM_INTERVALS-1) of integer;


--  function get_cdt_max_index (param      : integer) return integer;
--  function get_cdt_max_byte (param       : integer) return integer;
--  function get_cdt_max_byte_table (param : integer) return integer;
--  function get_reverse_table(param       : integer) return reverse_table_type;
--  function get_get_mul_factor(param      : integer) return integer;
--  function get_intervals_table(param     : integer) return intervals_type;
--  function get_intervals_table_max(param : integer) return intervals_type;


--end cdt_sampler_pkg;

--package body cdt_sampler_pkg is


--  function get_get_mul_factor(param : integer) return integer is
--  begin
--    if param = 1 then
--      return 8;
--    end if;
--  end get_get_mul_factor;


--  function get_cdt_max_byte_table (param : integer) return integer is
--  begin
--    if param = 1 then
--      return 9;
--    end if;
--  end get_cdt_max_byte_table;


--  function get_cdt_max_byte (param : integer) return integer is
--  begin
--    if param = 1 then
--      return 35;
--    end if;
--  end get_cdt_max_byte;


--  function get_cdt_max_index (param : integer) return integer is
--  begin
--    if param = 1 then
--      return 354;
--    end if;
--  end get_cdt_max_index;



--  function get_intervals_table(param : integer) return intervals_type is
--    constant intervals : intervals_type := (0, 353, 706, 1024, 1318, 1588, 1829, 2027, 2201, 2314, 0, 0, 0, 0, 0, 0);
--  begin
--    if param = 1 then
--      return intervals;
--    end if;
--  end get_intervals_table;


--  function get_intervals_table_max(param : integer) return intervals_type is
--    constant max_table : intervals_type := (353, 353, 318, 294, 270, 241, 198, 174, 113, 0, 0, 0, 0, 0, 0, 0);
--  begin
--    if param = 1 then
--      return max_table;
--    end if;
--  end get_intervals_table_max;


--  function get_reverse_table(param : integer) return reverse_table_type is
--    constant reverse_table_bliss_1 : reverse_table_type := ("1001101101100001", "1000111001001110", "1000011001001000", "1000000001000100", "0111110001000001", "0111100000111111", "0111011000111101", "0111001000111100", "0111000000111010", "0110111000111001", "0110110000111000", "0110101000110111", "0110100000110110", "0110011000110101", "0110010000110100", "0110010000110011", "0110001000110011", "0110000000110010", "0110000000110001", "0101111000110001", "0101110000110000", "0101110000101111", "0101101000101111", "0101101000101110", "0101100000101110", "0101100000101101", "0101011000101101", "0101011000101100", "0101010000101100", "0101010000101011", "0101001000101011", "0101001000101010", "0101000000101010", "0101000000101001", "0101000000101001", "0100111000101001", "0100111000101000", "0100111000101000", "0100110000101000", "0100110000100111", "0100101000100111", "0100101000100110", "0100101000100110", "0100100000100110", "0100100000100101", "0100100000100101", "0100011000100101", "0100011000100100", "0100011000100100", "0100011000100100", "0100010000100100", "0100010000100011", "0100010000100011", "0100001000100011", "0100001000100010", "0100001000100010", "0100001000100010", "0100000000100010", "0100000000100001", "0100000000100001", "0011111000100001", "0011111000100000", "0011111000100000", "0011111000100000", "0011110000100000", "0011110000011111", "0011110000011111", "0011110000011111", "0011101000011111", "0011101000011110", "0011101000011110", "0011101000011110", "0011101000011110", "0011100000011110", "0011100000011101", "0011100000011101", "0011100000011101", "0011011000011101", "0011011000011100", "0011011000011100", "0011011000011100", "0011011000011100", "0011010000011100", "0011010000011011", "0011010000011011", "0011010000011011", "0011001000011011", "0011001000011010", "0011001000011010", "0011001000011010", "0011001000011010", "0011000000011010", "0011000000011001", "0011000000011001", "0011000000011001", "0011000000011001", "0010111000011001", "0010111000011000", "0010111000011000", "0010111000011000", "0010111000011000", "0010111000011000", "0010110000011000", "0010110000010111", "0010110000010111", "0010110000010111", "0010110000010111", "0010101000010111", "0010101000010110", "0010101000010110", "0010101000010110", "0010101000010110", "0010101000010110", "0010100000010110", "0010100000010101", "0010100000010101", "0010100000010101", "0010100000010101", "0010011000010101", "0010011000010100", "0010011000010100", "0010011000010100", "0010011000010100", "0010011000010100", "0010010000010100", "0010010000010011", "0010010000010011", "0010010000010011", "0010010000010011", "0010010000010011", "0010001000010011", "0010001000010010", "0010001000010010", "0010001000010010", "0010001000010010", "0010001000010010", "0010001000010010", "0010000000010010", "0010000000010001", "0010000000010001", "0010000000010001", "0010000000010001", "0010000000010001", "0001111000010001", "0001111000010000", "0001111000010000", "0001111000010000", "0001111000010000", "0001111000010000", "0001111000010000", "0001110000010000", "0001110000001111", "0001110000001111", "0001110000001111", "0001110000001111", "0001110000001111", "0001101000001111", "0001101000001110", "0001101000001110", "0001101000001110", "0001101000001110", "0001101000001110", "0001101000001110", "0001100000001110", "0001100000001101", "0001100000001101", "0001100000001101", "0001100000001101", "0001100000001101", "0001100000001101", "0001011000001101", "0001011000001100", "0001011000001100", "0001011000001100", "0001011000001100", "0001011000001100", "0001011000001100", "0001010000001100", "0001010000001011", "0001010000001011", "0001010000001011", "0001010000001011", "0001010000001011", "0001010000001011", "0001001000001011", "0001001000001010", "0001001000001010", "0001001000001010", "0001001000001010", "0001001000001010", "0001001000001010", "0001000000001010", "0001000000001001", "0001000000001001", "0001000000001001", "0001000000001001", "0001000000001001", "0001000000001001", "0001000000001001", "0000111000001001", "0000111000001000", "0000111000001000", "0000111000001000", "0000111000001000", "0000111000001000", "0000111000001000", "0000110000001000", "0000110000000111", "0000110000000111", "0000110000000111", "0000110000000111", "0000110000000111", "0000110000000111", "0000110000000111", "0000101000000111", "0000101000000110", "0000101000000110", "0000101000000110", "0000101000000110", "0000101000000110", "0000101000000110", "0000100000000110", "0000100000000101", "0000100000000101", "0000100000000101", "0000100000000101", "0000100000000101", "0000100000000101", "0000100000000101", "0000011000000101", "0000011000000100", "0000011000000100", "0000011000000100", "0000011000000100", "0000011000000100", "0000011000000100", "0000010000000100", "0000010000000011", "0000010000000011", "0000010000000011", "0000010000000011", "0000010000000011", "0000010000000011", "0000010000000011", "0000001000000011", "0000001000000010", "0000001000000010", "0000001000000010", "0000001000000010", "0000001000000010", "0000001000000010", "0000001000000010", "0000000000000010", "0000000000000001", "0000000000000001", "0000000000000001");
--  begin
--    if param = 1 then
--      return reverse_table_bliss_1;
--    end if;
--  end get_reverse_table;



--end cdt_sampler_pkg;
